module BundleBridgeNexus_13(
  output  auto_out
);
  wire  outputs_0 = 1'h0; // @[HasTiles.scala 144:32]
  assign auto_out = outputs_0; // @[Nodes.scala 1213:84 BundleBridge.scala 151:67]
endmodule
