module IntSyncCrossingSource_1(
  input   auto_in_0,
  output  auto_out_sync_0
);
  assign auto_out_sync_0 = auto_in_0; // @[Nodes.scala 1216:84 LazyModule.scala 312:16]
endmodule
