module RVCExpander(
  input  [31:0] io_in,
  output [31:0] io_out_bits,
  output [4:0]  io_out_rd,
  output [4:0]  io_out_rs1,
  output [4:0]  io_out_rs2,
  output [4:0]  io_out_rs3,
  output        io_rvc
);
  wire [6:0] io_out_s_left_left = |(io_in[12:5]) ? 7'h13 : 7'h1f; // @[RVC.scala 54:20]
  wire [3:0] io_out_s_right_right_right = io_in[10:7]; // @[RVC.scala 35:26]
  wire [1:0] io_out_s_right_right_left = io_in[12:11]; // @[RVC.scala 35:35]
  wire  io_out_s_right_left = io_in[5]; // @[RVC.scala 35:45]
  wire  io_out_s_left_right = io_in[6]; // @[RVC.scala 35:51]
  wire [2:0] io_out_s_left_1 = io_in[4:2]; // @[RVC.scala 32:29]
  wire [4:0] io_out_s_left_right_1 = {2'h1,io_out_s_left_1}; // @[Cat.scala 29:58]
  wire [29:0] _io_out_s_T = {io_out_s_right_right_right,io_out_s_right_right_left,io_out_s_right_left,
    io_out_s_left_right,2'h0,5'h2,3'h0,2'h1,io_out_s_left_1,io_out_s_left_left}; // @[Cat.scala 29:58]
  wire [4:0] io_out_s_0_rs3 = io_in[31:27]; // @[RVC.scala 21:101]
  wire [1:0] io_out_s_right_right_2 = io_in[6:5]; // @[RVC.scala 37:20]
  wire [2:0] io_out_s_right_left_1 = io_in[12:10]; // @[RVC.scala 37:28]
  wire [7:0] io_out_s_right_right_right_2 = {io_out_s_right_right_2,io_out_s_right_left_1,3'h0}; // @[Cat.scala 29:58]
  wire [2:0] io_out_s_left_5 = io_in[9:7]; // @[RVC.scala 31:29]
  wire [4:0] io_out_s_right_right_left_1 = {2'h1,io_out_s_left_5}; // @[Cat.scala 29:58]
  wire [27:0] _io_out_s_T_4 = {io_out_s_right_right_2,io_out_s_right_left_1,3'h0,2'h1,io_out_s_left_5,3'h3,2'h1,
    io_out_s_left_1,7'h7}; // @[Cat.scala 29:58]
  wire [6:0] io_out_s_right_right_right_3 = {io_out_s_right_left,io_out_s_right_left_1,io_out_s_left_right,2'h0}; // @[Cat.scala 29:58]
  wire [26:0] _io_out_s_T_9 = {io_out_s_right_left,io_out_s_right_left_1,io_out_s_left_right,2'h0,2'h1,io_out_s_left_5,3'h2
    ,2'h1,io_out_s_left_1,7'h3}; // @[Cat.scala 29:58]
  wire [27:0] _io_out_s_T_14 = {io_out_s_right_right_2,io_out_s_right_left_1,3'h0,2'h1,io_out_s_left_5,3'h3,2'h1,
    io_out_s_left_1,7'h3}; // @[Cat.scala 29:58]
  wire [1:0] io_out_s_right_right_right_5 = io_out_s_right_right_right_3[6:5]; // @[RVC.scala 64:32]
  wire [4:0] io_out_s_left_right_left = io_out_s_right_right_right_3[4:0]; // @[RVC.scala 64:65]
  wire [26:0] _io_out_s_T_21 = {io_out_s_right_right_right_5,2'h1,io_out_s_left_1,2'h1,io_out_s_left_5,3'h2,
    io_out_s_left_right_left,7'h3f}; // @[Cat.scala 29:58]
  wire [2:0] io_out_s_right_right_right_6 = io_out_s_right_right_right_2[7:5]; // @[RVC.scala 67:30]
  wire [4:0] io_out_s_left_right_left_1 = io_out_s_right_right_right_2[4:0]; // @[RVC.scala 67:63]
  wire [27:0] _io_out_s_T_28 = {io_out_s_right_right_right_6,2'h1,io_out_s_left_1,2'h1,io_out_s_left_5,3'h3,
    io_out_s_left_right_left_1,7'h27}; // @[Cat.scala 29:58]
  wire [26:0] _io_out_s_T_35 = {io_out_s_right_right_right_5,2'h1,io_out_s_left_1,2'h1,io_out_s_left_5,3'h2,
    io_out_s_left_right_left,7'h23}; // @[Cat.scala 29:58]
  wire [27:0] _io_out_s_T_42 = {io_out_s_right_right_right_6,2'h1,io_out_s_left_1,2'h1,io_out_s_left_5,3'h3,
    io_out_s_left_right_left_1,7'h23}; // @[Cat.scala 29:58]
  wire [6:0] io_out_s_right_20 = io_in[12] ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12]
  wire [4:0] io_out_s_left_52 = io_in[6:2]; // @[RVC.scala 44:38]
  wire [11:0] io_out_s_right_right_right_9 = {io_out_s_right_20,io_out_s_left_52}; // @[Cat.scala 29:58]
  wire [4:0] io_out_s_right_right_left_8 = io_in[11:7]; // @[RVC.scala 34:13]
  wire [31:0] io_out_s_8_bits = {io_out_s_right_20,io_out_s_left_52,io_out_s_right_right_left_8,3'h0,
    io_out_s_right_right_left_8,7'h13}; // @[Cat.scala 29:58]
  wire  _io_out_s_opc_T_3 = |io_out_s_right_right_left_8; // @[RVC.scala 78:24]
  wire [6:0] io_out_s_left_left_1 = |io_out_s_right_right_left_8 ? 7'h1b : 7'h1f; // @[RVC.scala 78:20]
  wire [31:0] io_out_s_9_bits = {io_out_s_right_20,io_out_s_left_52,io_out_s_right_right_left_8,3'h0,
    io_out_s_right_right_left_8,io_out_s_left_left_1}; // @[Cat.scala 29:58]
  wire [31:0] io_out_s_10_bits = {io_out_s_right_20,io_out_s_left_52,5'h0,3'h0,io_out_s_right_right_left_8,7'h13}; // @[Cat.scala 29:58]
  wire  _io_out_s_opc_T_7 = |io_out_s_right_right_right_9; // @[RVC.scala 91:29]
  wire [6:0] io_out_s_me_left = |io_out_s_right_right_right_9 ? 7'h37 : 7'h3f; // @[RVC.scala 91:20]
  wire [14:0] io_out_s_me_right_right = io_in[12] ? 15'h7fff : 15'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _io_out_s_me_T_2 = {io_out_s_me_right_right,io_out_s_left_52,12'h0}; // @[Cat.scala 29:58]
  wire [19:0] io_out_s_me_right_right_1 = _io_out_s_me_T_2[31:12]; // @[RVC.scala 92:31]
  wire [31:0] io_out_s_me_bits = {io_out_s_me_right_right_1,io_out_s_right_right_left_8,io_out_s_me_left}; // @[Cat.scala 29:58]
  wire  _io_out_s_T_71 = (io_out_s_right_right_left_8 == 5'h0) | (io_out_s_right_right_left_8 == 5'h2); // @[RVC.scala 93:21]
  wire [6:0] io_out_s_left_left_2 = _io_out_s_opc_T_7 ? 7'h13 : 7'h1f; // @[RVC.scala 87:20]
  wire [2:0] io_out_s_right_right_right_12 = io_in[12] ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [1:0] io_out_s_right_right_left_10 = io_in[4:3]; // @[RVC.scala 43:42]
  wire  io_out_s_left_right_right = io_in[2]; // @[RVC.scala 43:56]
  wire [31:0] io_out_s_res_bits = {io_out_s_right_right_right_12,io_out_s_right_right_left_10,io_out_s_right_left,
    io_out_s_left_right_right,io_out_s_left_right,4'h0,io_out_s_right_right_left_8,3'h0,io_out_s_right_right_left_8,
    io_out_s_left_left_2}; // @[Cat.scala 29:58]
  wire [31:0] io_out_s_11_bits = _io_out_s_T_71 ? io_out_s_res_bits : io_out_s_me_bits; // @[RVC.scala 93:10]
  wire [4:0] io_out_s_11_rd = _io_out_s_T_71 ? io_out_s_right_right_left_8 : io_out_s_right_right_left_8; // @[RVC.scala 93:10]
  wire [4:0] io_out_s_11_rs2 = _io_out_s_T_71 ? io_out_s_left_right_1 : io_out_s_left_right_1; // @[RVC.scala 93:10]
  wire [4:0] io_out_s_11_rs3 = _io_out_s_T_71 ? io_out_s_0_rs3 : io_out_s_0_rs3; // @[RVC.scala 93:10]
  wire [25:0] _io_out_s_T_79 = {io_in[12],io_out_s_left_52,2'h1,io_out_s_left_5,3'h5,2'h1,io_out_s_left_5,7'h13}; // @[Cat.scala 29:58]
  wire [30:0] _GEN_0 = {{5'd0}, _io_out_s_T_79}; // @[RVC.scala 100:23]
  wire [30:0] _io_out_s_T_81 = _GEN_0 | 31'h40000000; // @[RVC.scala 100:23]
  wire [31:0] _io_out_s_T_84 = {io_out_s_right_20,io_out_s_left_52,2'h1,io_out_s_left_5,3'h7,2'h1,io_out_s_left_5,7'h13}
    ; // @[Cat.scala 29:58]
  wire [2:0] io_out_s_funct_truncIdx = {io_in[12],io_out_s_right_right_2}; // @[Cat.scala 29:58]
  wire [2:0] _io_out_s_funct_T_1 = io_out_s_funct_truncIdx == 3'h1 ? 3'h4 : 3'h0; // @[package.scala 32:76]
  wire [2:0] _io_out_s_funct_T_3 = io_out_s_funct_truncIdx == 3'h2 ? 3'h6 : _io_out_s_funct_T_1; // @[package.scala 32:76]
  wire [2:0] _io_out_s_funct_T_5 = io_out_s_funct_truncIdx == 3'h3 ? 3'h7 : _io_out_s_funct_T_3; // @[package.scala 32:76]
  wire [2:0] _io_out_s_funct_T_7 = io_out_s_funct_truncIdx == 3'h4 ? 3'h0 : _io_out_s_funct_T_5; // @[package.scala 32:76]
  wire [2:0] _io_out_s_funct_T_9 = io_out_s_funct_truncIdx == 3'h5 ? 3'h0 : _io_out_s_funct_T_7; // @[package.scala 32:76]
  wire [2:0] _io_out_s_funct_T_11 = io_out_s_funct_truncIdx == 3'h6 ? 3'h2 : _io_out_s_funct_T_9; // @[package.scala 32:76]
  wire [2:0] io_out_s_right_left_17 = io_out_s_funct_truncIdx == 3'h7 ? 3'h3 : _io_out_s_funct_T_11; // @[package.scala 32:76]
  wire [30:0] io_out_s_sub = io_out_s_right_right_2 == 2'h0 ? 31'h40000000 : 31'h0; // @[RVC.scala 104:22]
  wire [6:0] io_out_s_left_left_3 = io_in[12] ? 7'h3b : 7'h33; // @[RVC.scala 105:22]
  wire [24:0] _io_out_s_T_85 = {2'h1,io_out_s_left_1,2'h1,io_out_s_left_5,io_out_s_right_left_17,2'h1,io_out_s_left_5,
    io_out_s_left_left_3}; // @[Cat.scala 29:58]
  wire [30:0] _GEN_1 = {{6'd0}, _io_out_s_T_85}; // @[RVC.scala 106:43]
  wire [30:0] _io_out_s_T_86 = _GEN_1 | io_out_s_sub; // @[RVC.scala 106:43]
  wire [1:0] io_out_s_truncIdx = io_in[11:10]; // @[RVC.scala 108:42]
  wire [30:0] _io_out_s_T_88 = io_out_s_truncIdx == 2'h1 ? _io_out_s_T_81 : {{5'd0}, _io_out_s_T_79}; // @[package.scala 32:76]
  wire [31:0] _io_out_s_T_90 = io_out_s_truncIdx == 2'h2 ? _io_out_s_T_84 : {{1'd0}, _io_out_s_T_88}; // @[package.scala 32:76]
  wire [31:0] io_out_s_12_bits = io_out_s_truncIdx == 2'h3 ? {{1'd0}, _io_out_s_T_86} : _io_out_s_T_90; // @[package.scala 32:76]
  wire [9:0] io_out_s_right_right_right_right = io_in[12] ? 10'h3ff : 10'h0; // @[Bitwise.scala 72:12]
  wire  io_out_s_right_right_right_left = io_in[8]; // @[RVC.scala 45:36]
  wire [1:0] io_out_s_right_right_left_16 = io_in[10:9]; // @[RVC.scala 45:42]
  wire  io_out_s_right_left_left = io_in[7]; // @[RVC.scala 45:57]
  wire  io_out_s_left_right_left_5 = io_in[11]; // @[RVC.scala 45:69]
  wire [2:0] io_out_s_left_left_right = io_in[5:3]; // @[RVC.scala 45:76]
  wire [20:0] _io_out_s_T_99 = {io_out_s_right_right_right_right,io_out_s_right_right_right_left,
    io_out_s_right_right_left_16,io_out_s_left_right,io_out_s_right_left_left,io_out_s_left_right_right,
    io_out_s_left_right_left_5,io_out_s_left_left_right,1'h0}; // @[Cat.scala 29:58]
  wire  io_out_s_right_right_right_19 = _io_out_s_T_99[20]; // @[RVC.scala 95:26]
  wire [9:0] io_out_s_right_right_left_18 = _io_out_s_T_99[10:1]; // @[RVC.scala 95:36]
  wire  io_out_s_right_left_21 = _io_out_s_T_99[11]; // @[RVC.scala 95:48]
  wire [7:0] io_out_s_left_right_right_5 = _io_out_s_T_99[19:12]; // @[RVC.scala 95:58]
  wire [31:0] io_out_s_13_bits = {io_out_s_right_right_right_19,io_out_s_right_right_left_18,io_out_s_right_left_21,
    io_out_s_left_right_right_5,5'h0,7'h6f}; // @[Cat.scala 29:58]
  wire [4:0] io_out_s_right_right_right_23 = io_in[12] ? 5'h1f : 5'h0; // @[Bitwise.scala 72:12]
  wire [12:0] _io_out_s_T_115 = {io_out_s_right_right_right_23,io_out_s_right_right_2,io_out_s_left_right_right,
    io_out_s_truncIdx,io_out_s_right_right_left_10,1'h0}; // @[Cat.scala 29:58]
  wire  io_out_s_right_right_right_24 = _io_out_s_T_115[12]; // @[RVC.scala 96:29]
  wire [5:0] io_out_s_right_right_left_23 = _io_out_s_T_115[10:5]; // @[RVC.scala 96:39]
  wire [3:0] io_out_s_left_right_left_12 = _io_out_s_T_115[4:1]; // @[RVC.scala 96:71]
  wire  io_out_s_left_left_right_4 = _io_out_s_T_115[11]; // @[RVC.scala 96:82]
  wire [31:0] io_out_s_14_bits = {io_out_s_right_right_right_24,io_out_s_right_right_left_23,5'h0,2'h1,io_out_s_left_5,3'h0
    ,io_out_s_left_right_left_12,io_out_s_left_left_right_4,7'h63}; // @[Cat.scala 29:58]
  wire [31:0] io_out_s_15_bits = {io_out_s_right_right_right_24,io_out_s_right_right_left_23,5'h0,2'h1,io_out_s_left_5,3'h1
    ,io_out_s_left_right_left_12,io_out_s_left_left_right_4,7'h63}; // @[Cat.scala 29:58]
  wire [6:0] io_out_s_left_left_10 = _io_out_s_opc_T_3 ? 7'h3 : 7'h1f; // @[RVC.scala 114:23]
  wire [25:0] _io_out_s_T_144 = {io_in[12],io_out_s_left_52,io_out_s_right_right_left_8,3'h1,io_out_s_right_right_left_8
    ,7'h13}; // @[Cat.scala 29:58]
  wire [28:0] _io_out_s_T_149 = {io_out_s_left_1,io_in[12],io_out_s_right_right_2,3'h0,5'h2,3'h3,
    io_out_s_right_right_left_8,7'h7}; // @[Cat.scala 29:58]
  wire [1:0] io_out_s_right_right_47 = io_in[3:2]; // @[RVC.scala 38:22]
  wire [2:0] io_out_s_left_right_41 = io_in[6:4]; // @[RVC.scala 38:37]
  wire [27:0] _io_out_s_T_153 = {io_out_s_right_right_47,io_in[12],io_out_s_left_right_41,2'h0,5'h2,3'h2,
    io_out_s_right_right_left_8,io_out_s_left_left_10}; // @[Cat.scala 29:58]
  wire [28:0] _io_out_s_T_157 = {io_out_s_left_1,io_in[12],io_out_s_right_right_2,3'h0,5'h2,3'h3,
    io_out_s_right_right_left_8,io_out_s_left_left_10}; // @[Cat.scala 29:58]
  wire [24:0] _io_out_s_mv_T = {io_out_s_left_52,5'h0,3'h0,io_out_s_right_right_left_8,7'h33}; // @[Cat.scala 29:58]
  wire [24:0] _io_out_s_add_T = {io_out_s_left_52,io_out_s_right_right_left_8,3'h0,io_out_s_right_right_left_8,7'h33}; // @[Cat.scala 29:58]
  wire [24:0] io_out_s_jr = {io_out_s_left_52,io_out_s_right_right_left_8,3'h0,12'h67}; // @[Cat.scala 29:58]
  wire [17:0] io_out_s_reserved_right = io_out_s_jr[24:7]; // @[RVC.scala 134:29]
  wire [24:0] io_out_s_reserved = {io_out_s_reserved_right,7'h1f}; // @[Cat.scala 29:58]
  wire [24:0] _io_out_s_jr_reserved_T_2 = _io_out_s_opc_T_3 ? io_out_s_jr : io_out_s_reserved; // @[RVC.scala 135:33]
  wire  _io_out_s_jr_mv_T_1 = |io_out_s_left_52; // @[RVC.scala 136:27]
  wire [31:0] io_out_s_mv_bits = {{7'd0}, _io_out_s_mv_T}; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] io_out_s_jr_reserved_bits = {{7'd0}, _io_out_s_jr_reserved_T_2}; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] io_out_s_jr_mv_bits = |io_out_s_left_52 ? io_out_s_mv_bits : io_out_s_jr_reserved_bits; // @[RVC.scala 136:22]
  wire [4:0] io_out_s_jr_mv_rd = |io_out_s_left_52 ? io_out_s_right_right_left_8 : 5'h0; // @[RVC.scala 136:22]
  wire [4:0] io_out_s_jr_mv_rs1 = |io_out_s_left_52 ? 5'h0 : io_out_s_right_right_left_8; // @[RVC.scala 136:22]
  wire [4:0] io_out_s_jr_mv_rs2 = |io_out_s_left_52 ? io_out_s_left_52 : io_out_s_left_52; // @[RVC.scala 136:22]
  wire [4:0] io_out_s_jr_mv_rs3 = |io_out_s_left_52 ? io_out_s_0_rs3 : io_out_s_0_rs3; // @[RVC.scala 136:22]
  wire [24:0] io_out_s_jalr = {io_out_s_left_52,io_out_s_right_right_left_8,3'h0,12'he7}; // @[Cat.scala 29:58]
  wire [24:0] _io_out_s_ebreak_T = {io_out_s_reserved_right,7'h73}; // @[Cat.scala 29:58]
  wire [24:0] io_out_s_ebreak = _io_out_s_ebreak_T | 25'h100000; // @[RVC.scala 138:46]
  wire [24:0] _io_out_s_jalr_ebreak_T_2 = _io_out_s_opc_T_3 ? io_out_s_jalr : io_out_s_ebreak; // @[RVC.scala 139:33]
  wire [31:0] io_out_s_add_bits = {{7'd0}, _io_out_s_add_T}; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] io_out_s_jalr_ebreak_bits = {{7'd0}, _io_out_s_jalr_ebreak_T_2}; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] io_out_s_jalr_add_bits = _io_out_s_jr_mv_T_1 ? io_out_s_add_bits : io_out_s_jalr_ebreak_bits; // @[RVC.scala 140:25]
  wire [4:0] io_out_s_jalr_add_rd = _io_out_s_jr_mv_T_1 ? io_out_s_right_right_left_8 : 5'h1; // @[RVC.scala 140:25]
  wire [4:0] io_out_s_jalr_add_rs1 = _io_out_s_jr_mv_T_1 ? io_out_s_right_right_left_8 : io_out_s_right_right_left_8; // @[RVC.scala 140:25]
  wire [31:0] io_out_s_20_bits = io_in[12] ? io_out_s_jalr_add_bits : io_out_s_jr_mv_bits; // @[RVC.scala 141:10]
  wire [4:0] io_out_s_20_rd = io_in[12] ? io_out_s_jalr_add_rd : io_out_s_jr_mv_rd; // @[RVC.scala 141:10]
  wire [4:0] io_out_s_20_rs1 = io_in[12] ? io_out_s_jalr_add_rs1 : io_out_s_jr_mv_rs1; // @[RVC.scala 141:10]
  wire [4:0] io_out_s_20_rs2 = io_in[12] ? io_out_s_jr_mv_rs2 : io_out_s_jr_mv_rs2; // @[RVC.scala 141:10]
  wire [4:0] io_out_s_20_rs3 = io_in[12] ? io_out_s_jr_mv_rs3 : io_out_s_jr_mv_rs3; // @[RVC.scala 141:10]
  wire [8:0] _io_out_s_T_162 = {io_out_s_left_5,io_out_s_right_left_1,3'h0}; // @[Cat.scala 29:58]
  wire [3:0] io_out_s_right_right_right_37 = _io_out_s_T_162[8:5]; // @[RVC.scala 125:34]
  wire [4:0] io_out_s_left_right_left_19 = _io_out_s_T_162[4:0]; // @[RVC.scala 125:66]
  wire [28:0] _io_out_s_T_164 = {io_out_s_right_right_right_37,io_out_s_left_52,5'h2,3'h3,io_out_s_left_right_left_19,7'h27
    }; // @[Cat.scala 29:58]
  wire [1:0] io_out_s_right_right_54 = io_in[8:7]; // @[RVC.scala 40:22]
  wire [3:0] io_out_s_right_left_38 = io_in[12:9]; // @[RVC.scala 40:30]
  wire [7:0] _io_out_s_T_168 = {io_out_s_right_right_54,io_out_s_right_left_38,2'h0}; // @[Cat.scala 29:58]
  wire [2:0] io_out_s_right_right_right_38 = _io_out_s_T_168[7:5]; // @[RVC.scala 124:33]
  wire [4:0] io_out_s_left_right_left_20 = _io_out_s_T_168[4:0]; // @[RVC.scala 124:65]
  wire [27:0] _io_out_s_T_170 = {io_out_s_right_right_right_38,io_out_s_left_52,5'h2,3'h2,io_out_s_left_right_left_20,7'h23
    }; // @[Cat.scala 29:58]
  wire [28:0] _io_out_s_T_176 = {io_out_s_right_right_right_37,io_out_s_left_52,5'h2,3'h3,io_out_s_left_right_left_19,7'h23
    }; // @[Cat.scala 29:58]
  wire [4:0] io_out_s_24_rs1 = io_in[19:15]; // @[RVC.scala 21:57]
  wire [4:0] io_out_s_24_rs2 = io_in[24:20]; // @[RVC.scala 21:79]
  wire [2:0] io_out_left = io_in[15:13]; // @[RVC.scala 152:20]
  wire [4:0] io_out_truncIdx = {io_in[1:0],io_out_left}; // @[Cat.scala 29:58]
  wire [31:0] io_out_s_1_bits = {{4'd0}, _io_out_s_T_4}; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] io_out_s_0_bits = {{2'd0}, _io_out_s_T}; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] _io_out_T_1_bits = io_out_truncIdx == 5'h1 ? io_out_s_1_bits : io_out_s_0_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_1_rd = io_out_truncIdx == 5'h1 ? io_out_s_left_right_1 : io_out_s_left_right_1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_1_rs1 = io_out_truncIdx == 5'h1 ? io_out_s_right_right_left_1 : 5'h2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_1_rs3 = io_out_truncIdx == 5'h1 ? io_out_s_0_rs3 : io_out_s_0_rs3; // @[package.scala 32:76]
  wire [31:0] io_out_s_2_bits = {{5'd0}, _io_out_s_T_9}; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] _io_out_T_3_bits = io_out_truncIdx == 5'h2 ? io_out_s_2_bits : _io_out_T_1_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_3_rd = io_out_truncIdx == 5'h2 ? io_out_s_left_right_1 : _io_out_T_1_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_3_rs1 = io_out_truncIdx == 5'h2 ? io_out_s_right_right_left_1 : _io_out_T_1_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_3_rs3 = io_out_truncIdx == 5'h2 ? io_out_s_0_rs3 : _io_out_T_1_rs3; // @[package.scala 32:76]
  wire [31:0] io_out_s_3_bits = {{4'd0}, _io_out_s_T_14}; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] _io_out_T_5_bits = io_out_truncIdx == 5'h3 ? io_out_s_3_bits : _io_out_T_3_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_5_rd = io_out_truncIdx == 5'h3 ? io_out_s_left_right_1 : _io_out_T_3_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_5_rs1 = io_out_truncIdx == 5'h3 ? io_out_s_right_right_left_1 : _io_out_T_3_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_5_rs3 = io_out_truncIdx == 5'h3 ? io_out_s_0_rs3 : _io_out_T_3_rs3; // @[package.scala 32:76]
  wire [31:0] io_out_s_4_bits = {{5'd0}, _io_out_s_T_21}; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] _io_out_T_7_bits = io_out_truncIdx == 5'h4 ? io_out_s_4_bits : _io_out_T_5_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_7_rd = io_out_truncIdx == 5'h4 ? io_out_s_left_right_1 : _io_out_T_5_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_7_rs1 = io_out_truncIdx == 5'h4 ? io_out_s_right_right_left_1 : _io_out_T_5_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_7_rs3 = io_out_truncIdx == 5'h4 ? io_out_s_0_rs3 : _io_out_T_5_rs3; // @[package.scala 32:76]
  wire [31:0] io_out_s_5_bits = {{4'd0}, _io_out_s_T_28}; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] _io_out_T_9_bits = io_out_truncIdx == 5'h5 ? io_out_s_5_bits : _io_out_T_7_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_9_rd = io_out_truncIdx == 5'h5 ? io_out_s_left_right_1 : _io_out_T_7_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_9_rs1 = io_out_truncIdx == 5'h5 ? io_out_s_right_right_left_1 : _io_out_T_7_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_9_rs3 = io_out_truncIdx == 5'h5 ? io_out_s_0_rs3 : _io_out_T_7_rs3; // @[package.scala 32:76]
  wire [31:0] io_out_s_6_bits = {{5'd0}, _io_out_s_T_35}; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] _io_out_T_11_bits = io_out_truncIdx == 5'h6 ? io_out_s_6_bits : _io_out_T_9_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_11_rd = io_out_truncIdx == 5'h6 ? io_out_s_left_right_1 : _io_out_T_9_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_11_rs1 = io_out_truncIdx == 5'h6 ? io_out_s_right_right_left_1 : _io_out_T_9_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_11_rs3 = io_out_truncIdx == 5'h6 ? io_out_s_0_rs3 : _io_out_T_9_rs3; // @[package.scala 32:76]
  wire [31:0] io_out_s_7_bits = {{4'd0}, _io_out_s_T_42}; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] _io_out_T_13_bits = io_out_truncIdx == 5'h7 ? io_out_s_7_bits : _io_out_T_11_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_13_rd = io_out_truncIdx == 5'h7 ? io_out_s_left_right_1 : _io_out_T_11_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_13_rs1 = io_out_truncIdx == 5'h7 ? io_out_s_right_right_left_1 : _io_out_T_11_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_13_rs3 = io_out_truncIdx == 5'h7 ? io_out_s_0_rs3 : _io_out_T_11_rs3; // @[package.scala 32:76]
  wire [31:0] _io_out_T_15_bits = io_out_truncIdx == 5'h8 ? io_out_s_8_bits : _io_out_T_13_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_15_rd = io_out_truncIdx == 5'h8 ? io_out_s_right_right_left_8 : _io_out_T_13_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_15_rs1 = io_out_truncIdx == 5'h8 ? io_out_s_right_right_left_8 : _io_out_T_13_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_15_rs2 = io_out_truncIdx == 5'h8 ? io_out_s_left_right_1 : _io_out_T_13_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_15_rs3 = io_out_truncIdx == 5'h8 ? io_out_s_0_rs3 : _io_out_T_13_rs3; // @[package.scala 32:76]
  wire [31:0] _io_out_T_17_bits = io_out_truncIdx == 5'h9 ? io_out_s_9_bits : _io_out_T_15_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_17_rd = io_out_truncIdx == 5'h9 ? io_out_s_right_right_left_8 : _io_out_T_15_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_17_rs1 = io_out_truncIdx == 5'h9 ? io_out_s_right_right_left_8 : _io_out_T_15_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_17_rs2 = io_out_truncIdx == 5'h9 ? io_out_s_left_right_1 : _io_out_T_15_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_17_rs3 = io_out_truncIdx == 5'h9 ? io_out_s_0_rs3 : _io_out_T_15_rs3; // @[package.scala 32:76]
  wire [31:0] _io_out_T_19_bits = io_out_truncIdx == 5'ha ? io_out_s_10_bits : _io_out_T_17_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_19_rd = io_out_truncIdx == 5'ha ? io_out_s_right_right_left_8 : _io_out_T_17_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_19_rs1 = io_out_truncIdx == 5'ha ? 5'h0 : _io_out_T_17_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_19_rs2 = io_out_truncIdx == 5'ha ? io_out_s_left_right_1 : _io_out_T_17_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_19_rs3 = io_out_truncIdx == 5'ha ? io_out_s_0_rs3 : _io_out_T_17_rs3; // @[package.scala 32:76]
  wire [31:0] _io_out_T_21_bits = io_out_truncIdx == 5'hb ? io_out_s_11_bits : _io_out_T_19_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_21_rd = io_out_truncIdx == 5'hb ? io_out_s_11_rd : _io_out_T_19_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_21_rs1 = io_out_truncIdx == 5'hb ? io_out_s_11_rd : _io_out_T_19_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_21_rs2 = io_out_truncIdx == 5'hb ? io_out_s_11_rs2 : _io_out_T_19_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_21_rs3 = io_out_truncIdx == 5'hb ? io_out_s_11_rs3 : _io_out_T_19_rs3; // @[package.scala 32:76]
  wire [31:0] _io_out_T_23_bits = io_out_truncIdx == 5'hc ? io_out_s_12_bits : _io_out_T_21_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_23_rd = io_out_truncIdx == 5'hc ? io_out_s_right_right_left_1 : _io_out_T_21_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_23_rs1 = io_out_truncIdx == 5'hc ? io_out_s_right_right_left_1 : _io_out_T_21_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_23_rs2 = io_out_truncIdx == 5'hc ? io_out_s_left_right_1 : _io_out_T_21_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_23_rs3 = io_out_truncIdx == 5'hc ? io_out_s_0_rs3 : _io_out_T_21_rs3; // @[package.scala 32:76]
  wire [31:0] _io_out_T_25_bits = io_out_truncIdx == 5'hd ? io_out_s_13_bits : _io_out_T_23_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_25_rd = io_out_truncIdx == 5'hd ? 5'h0 : _io_out_T_23_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_25_rs1 = io_out_truncIdx == 5'hd ? io_out_s_right_right_left_1 : _io_out_T_23_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_25_rs2 = io_out_truncIdx == 5'hd ? io_out_s_left_right_1 : _io_out_T_23_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_25_rs3 = io_out_truncIdx == 5'hd ? io_out_s_0_rs3 : _io_out_T_23_rs3; // @[package.scala 32:76]
  wire [31:0] _io_out_T_27_bits = io_out_truncIdx == 5'he ? io_out_s_14_bits : _io_out_T_25_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_27_rd = io_out_truncIdx == 5'he ? io_out_s_right_right_left_1 : _io_out_T_25_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_27_rs1 = io_out_truncIdx == 5'he ? io_out_s_right_right_left_1 : _io_out_T_25_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_27_rs2 = io_out_truncIdx == 5'he ? 5'h0 : _io_out_T_25_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_27_rs3 = io_out_truncIdx == 5'he ? io_out_s_0_rs3 : _io_out_T_25_rs3; // @[package.scala 32:76]
  wire [31:0] _io_out_T_29_bits = io_out_truncIdx == 5'hf ? io_out_s_15_bits : _io_out_T_27_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_29_rd = io_out_truncIdx == 5'hf ? 5'h0 : _io_out_T_27_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_29_rs1 = io_out_truncIdx == 5'hf ? io_out_s_right_right_left_1 : _io_out_T_27_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_29_rs2 = io_out_truncIdx == 5'hf ? 5'h0 : _io_out_T_27_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_29_rs3 = io_out_truncIdx == 5'hf ? io_out_s_0_rs3 : _io_out_T_27_rs3; // @[package.scala 32:76]
  wire [31:0] io_out_s_16_bits = {{6'd0}, _io_out_s_T_144}; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] _io_out_T_31_bits = io_out_truncIdx == 5'h10 ? io_out_s_16_bits : _io_out_T_29_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_31_rd = io_out_truncIdx == 5'h10 ? io_out_s_right_right_left_8 : _io_out_T_29_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_31_rs1 = io_out_truncIdx == 5'h10 ? io_out_s_right_right_left_8 : _io_out_T_29_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_31_rs2 = io_out_truncIdx == 5'h10 ? io_out_s_left_52 : _io_out_T_29_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_31_rs3 = io_out_truncIdx == 5'h10 ? io_out_s_0_rs3 : _io_out_T_29_rs3; // @[package.scala 32:76]
  wire [31:0] io_out_s_17_bits = {{3'd0}, _io_out_s_T_149}; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] _io_out_T_33_bits = io_out_truncIdx == 5'h11 ? io_out_s_17_bits : _io_out_T_31_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_33_rd = io_out_truncIdx == 5'h11 ? io_out_s_right_right_left_8 : _io_out_T_31_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_33_rs1 = io_out_truncIdx == 5'h11 ? 5'h2 : _io_out_T_31_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_33_rs2 = io_out_truncIdx == 5'h11 ? io_out_s_left_52 : _io_out_T_31_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_33_rs3 = io_out_truncIdx == 5'h11 ? io_out_s_0_rs3 : _io_out_T_31_rs3; // @[package.scala 32:76]
  wire [31:0] io_out_s_18_bits = {{4'd0}, _io_out_s_T_153}; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] _io_out_T_35_bits = io_out_truncIdx == 5'h12 ? io_out_s_18_bits : _io_out_T_33_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_35_rd = io_out_truncIdx == 5'h12 ? io_out_s_right_right_left_8 : _io_out_T_33_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_35_rs1 = io_out_truncIdx == 5'h12 ? 5'h2 : _io_out_T_33_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_35_rs2 = io_out_truncIdx == 5'h12 ? io_out_s_left_52 : _io_out_T_33_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_35_rs3 = io_out_truncIdx == 5'h12 ? io_out_s_0_rs3 : _io_out_T_33_rs3; // @[package.scala 32:76]
  wire [31:0] io_out_s_19_bits = {{3'd0}, _io_out_s_T_157}; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] _io_out_T_37_bits = io_out_truncIdx == 5'h13 ? io_out_s_19_bits : _io_out_T_35_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_37_rd = io_out_truncIdx == 5'h13 ? io_out_s_right_right_left_8 : _io_out_T_35_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_37_rs1 = io_out_truncIdx == 5'h13 ? 5'h2 : _io_out_T_35_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_37_rs2 = io_out_truncIdx == 5'h13 ? io_out_s_left_52 : _io_out_T_35_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_37_rs3 = io_out_truncIdx == 5'h13 ? io_out_s_0_rs3 : _io_out_T_35_rs3; // @[package.scala 32:76]
  wire [31:0] _io_out_T_39_bits = io_out_truncIdx == 5'h14 ? io_out_s_20_bits : _io_out_T_37_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_39_rd = io_out_truncIdx == 5'h14 ? io_out_s_20_rd : _io_out_T_37_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_39_rs1 = io_out_truncIdx == 5'h14 ? io_out_s_20_rs1 : _io_out_T_37_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_39_rs2 = io_out_truncIdx == 5'h14 ? io_out_s_20_rs2 : _io_out_T_37_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_39_rs3 = io_out_truncIdx == 5'h14 ? io_out_s_20_rs3 : _io_out_T_37_rs3; // @[package.scala 32:76]
  wire [31:0] io_out_s_21_bits = {{3'd0}, _io_out_s_T_164}; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] _io_out_T_41_bits = io_out_truncIdx == 5'h15 ? io_out_s_21_bits : _io_out_T_39_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_41_rd = io_out_truncIdx == 5'h15 ? io_out_s_right_right_left_8 : _io_out_T_39_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_41_rs1 = io_out_truncIdx == 5'h15 ? 5'h2 : _io_out_T_39_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_41_rs2 = io_out_truncIdx == 5'h15 ? io_out_s_left_52 : _io_out_T_39_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_41_rs3 = io_out_truncIdx == 5'h15 ? io_out_s_0_rs3 : _io_out_T_39_rs3; // @[package.scala 32:76]
  wire [31:0] io_out_s_22_bits = {{4'd0}, _io_out_s_T_170}; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] _io_out_T_43_bits = io_out_truncIdx == 5'h16 ? io_out_s_22_bits : _io_out_T_41_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_43_rd = io_out_truncIdx == 5'h16 ? io_out_s_right_right_left_8 : _io_out_T_41_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_43_rs1 = io_out_truncIdx == 5'h16 ? 5'h2 : _io_out_T_41_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_43_rs2 = io_out_truncIdx == 5'h16 ? io_out_s_left_52 : _io_out_T_41_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_43_rs3 = io_out_truncIdx == 5'h16 ? io_out_s_0_rs3 : _io_out_T_41_rs3; // @[package.scala 32:76]
  wire [31:0] io_out_s_23_bits = {{3'd0}, _io_out_s_T_176}; // @[RVC.scala 22:19 RVC.scala 23:14]
  wire [31:0] _io_out_T_45_bits = io_out_truncIdx == 5'h17 ? io_out_s_23_bits : _io_out_T_43_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_45_rd = io_out_truncIdx == 5'h17 ? io_out_s_right_right_left_8 : _io_out_T_43_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_45_rs1 = io_out_truncIdx == 5'h17 ? 5'h2 : _io_out_T_43_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_45_rs2 = io_out_truncIdx == 5'h17 ? io_out_s_left_52 : _io_out_T_43_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_45_rs3 = io_out_truncIdx == 5'h17 ? io_out_s_0_rs3 : _io_out_T_43_rs3; // @[package.scala 32:76]
  wire [31:0] _io_out_T_47_bits = io_out_truncIdx == 5'h18 ? io_in : _io_out_T_45_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_47_rd = io_out_truncIdx == 5'h18 ? io_out_s_right_right_left_8 : _io_out_T_45_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_47_rs1 = io_out_truncIdx == 5'h18 ? io_out_s_24_rs1 : _io_out_T_45_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_47_rs2 = io_out_truncIdx == 5'h18 ? io_out_s_24_rs2 : _io_out_T_45_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_47_rs3 = io_out_truncIdx == 5'h18 ? io_out_s_0_rs3 : _io_out_T_45_rs3; // @[package.scala 32:76]
  wire [31:0] _io_out_T_49_bits = io_out_truncIdx == 5'h19 ? io_in : _io_out_T_47_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_49_rd = io_out_truncIdx == 5'h19 ? io_out_s_right_right_left_8 : _io_out_T_47_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_49_rs1 = io_out_truncIdx == 5'h19 ? io_out_s_24_rs1 : _io_out_T_47_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_49_rs2 = io_out_truncIdx == 5'h19 ? io_out_s_24_rs2 : _io_out_T_47_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_49_rs3 = io_out_truncIdx == 5'h19 ? io_out_s_0_rs3 : _io_out_T_47_rs3; // @[package.scala 32:76]
  wire [31:0] _io_out_T_51_bits = io_out_truncIdx == 5'h1a ? io_in : _io_out_T_49_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_51_rd = io_out_truncIdx == 5'h1a ? io_out_s_right_right_left_8 : _io_out_T_49_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_51_rs1 = io_out_truncIdx == 5'h1a ? io_out_s_24_rs1 : _io_out_T_49_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_51_rs2 = io_out_truncIdx == 5'h1a ? io_out_s_24_rs2 : _io_out_T_49_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_51_rs3 = io_out_truncIdx == 5'h1a ? io_out_s_0_rs3 : _io_out_T_49_rs3; // @[package.scala 32:76]
  wire [31:0] _io_out_T_53_bits = io_out_truncIdx == 5'h1b ? io_in : _io_out_T_51_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_53_rd = io_out_truncIdx == 5'h1b ? io_out_s_right_right_left_8 : _io_out_T_51_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_53_rs1 = io_out_truncIdx == 5'h1b ? io_out_s_24_rs1 : _io_out_T_51_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_53_rs2 = io_out_truncIdx == 5'h1b ? io_out_s_24_rs2 : _io_out_T_51_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_53_rs3 = io_out_truncIdx == 5'h1b ? io_out_s_0_rs3 : _io_out_T_51_rs3; // @[package.scala 32:76]
  wire [31:0] _io_out_T_55_bits = io_out_truncIdx == 5'h1c ? io_in : _io_out_T_53_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_55_rd = io_out_truncIdx == 5'h1c ? io_out_s_right_right_left_8 : _io_out_T_53_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_55_rs1 = io_out_truncIdx == 5'h1c ? io_out_s_24_rs1 : _io_out_T_53_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_55_rs2 = io_out_truncIdx == 5'h1c ? io_out_s_24_rs2 : _io_out_T_53_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_55_rs3 = io_out_truncIdx == 5'h1c ? io_out_s_0_rs3 : _io_out_T_53_rs3; // @[package.scala 32:76]
  wire [31:0] _io_out_T_57_bits = io_out_truncIdx == 5'h1d ? io_in : _io_out_T_55_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_57_rd = io_out_truncIdx == 5'h1d ? io_out_s_right_right_left_8 : _io_out_T_55_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_57_rs1 = io_out_truncIdx == 5'h1d ? io_out_s_24_rs1 : _io_out_T_55_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_57_rs2 = io_out_truncIdx == 5'h1d ? io_out_s_24_rs2 : _io_out_T_55_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_57_rs3 = io_out_truncIdx == 5'h1d ? io_out_s_0_rs3 : _io_out_T_55_rs3; // @[package.scala 32:76]
  wire [31:0] _io_out_T_59_bits = io_out_truncIdx == 5'h1e ? io_in : _io_out_T_57_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_59_rd = io_out_truncIdx == 5'h1e ? io_out_s_right_right_left_8 : _io_out_T_57_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_59_rs1 = io_out_truncIdx == 5'h1e ? io_out_s_24_rs1 : _io_out_T_57_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_59_rs2 = io_out_truncIdx == 5'h1e ? io_out_s_24_rs2 : _io_out_T_57_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_59_rs3 = io_out_truncIdx == 5'h1e ? io_out_s_0_rs3 : _io_out_T_57_rs3; // @[package.scala 32:76]
  assign io_out_bits = io_out_truncIdx == 5'h1f ? io_in : _io_out_T_59_bits; // @[package.scala 32:76]
  assign io_out_rd = io_out_truncIdx == 5'h1f ? io_out_s_right_right_left_8 : _io_out_T_59_rd; // @[package.scala 32:76]
  assign io_out_rs1 = io_out_truncIdx == 5'h1f ? io_out_s_24_rs1 : _io_out_T_59_rs1; // @[package.scala 32:76]
  assign io_out_rs2 = io_out_truncIdx == 5'h1f ? io_out_s_24_rs2 : _io_out_T_59_rs2; // @[package.scala 32:76]
  assign io_out_rs3 = io_out_truncIdx == 5'h1f ? io_out_s_0_rs3 : _io_out_T_59_rs3; // @[package.scala 32:76]
  assign io_rvc = (io_in[1:0]) != 2'h3; // @[RVC.scala 164:26]
endmodule
