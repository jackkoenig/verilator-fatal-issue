module OptimizationBarrier_117(
  input  [2:0] io_x,
  output [2:0] io_y
);
  assign io_y = io_x; // @[package.scala 241:12]
endmodule
