module RoundAnyRawFNToRecFN_3(
  input         io_invalidExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [12:0] io_in_sExp,
  input  [53:0] io_in_sig,
  input  [2:0]  io_roundingMode,
  output [32:0] io_out,
  output [4:0]  io_exceptionFlags
);
  wire  roundingMode_near_even = io_roundingMode == 3'h0; // @[RoundAnyRawFNToRecFN.scala 88:53]
  wire  roundingMode_min = io_roundingMode == 3'h2; // @[RoundAnyRawFNToRecFN.scala 90:53]
  wire  roundingMode_max = io_roundingMode == 3'h3; // @[RoundAnyRawFNToRecFN.scala 91:53]
  wire  roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RoundAnyRawFNToRecFN.scala 92:53]
  wire  roundingMode_odd = io_roundingMode == 3'h6; // @[RoundAnyRawFNToRecFN.scala 93:53]
  wire  roundMagUp = (roundingMode_min & io_in_sign) | (roundingMode_max & (~io_in_sign)); // @[RoundAnyRawFNToRecFN.scala 96:42]
  wire [13:0] sAdjustedExp = $signed(io_in_sExp) - 13'sh700; // @[RoundAnyRawFNToRecFN.scala 108:24]
  wire [25:0] adjustedSig_right = io_in_sig[53:28]; // @[RoundAnyRawFNToRecFN.scala 114:26]
  wire  adjustedSig_left = |(io_in_sig[27:0]); // @[RoundAnyRawFNToRecFN.scala 115:60]
  wire [26:0] adjustedSig = {adjustedSig_right,adjustedSig_left}; // @[Cat.scala 29:58]
  wire [8:0] _roundMask_T_1 = ~(sAdjustedExp[8:0]); // @[primitives.scala 51:21]
  wire  roundMask_msb = _roundMask_T_1[8]; // @[primitives.scala 57:25]
  wire [7:0] roundMask_lsbs = _roundMask_T_1[7:0]; // @[primitives.scala 58:26]
  wire  roundMask_msb_1 = roundMask_lsbs[7]; // @[primitives.scala 57:25]
  wire [6:0] roundMask_lsbs_1 = roundMask_lsbs[6:0]; // @[primitives.scala 58:26]
  wire  roundMask_msb_2 = roundMask_lsbs_1[6]; // @[primitives.scala 57:25]
  wire [5:0] roundMask_lsbs_2 = roundMask_lsbs_1[5:0]; // @[primitives.scala 58:26]
  wire [64:0] roundMask_shift = -65'sh10000000000000000 >>> roundMask_lsbs_2; // @[primitives.scala 77:58]
  wire [15:0] roundMask_res = roundMask_shift[57:42]; // @[Bitwise.scala 109:18]
  wire [15:0] _roundMask_T_6 = {{8'd0}, roundMask_res[15:8]}; // @[Bitwise.scala 103:31]
  wire [15:0] _roundMask_T_8 = {roundMask_res[7:0], 8'h0}; // @[Bitwise.scala 103:65]
  wire [15:0] _roundMask_T_10 = _roundMask_T_8 & 16'hff00; // @[Bitwise.scala 103:75]
  wire [15:0] _roundMask_T_11 = _roundMask_T_6 | _roundMask_T_10; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_0 = {{4'd0}, _roundMask_T_11[15:4]}; // @[Bitwise.scala 103:31]
  wire [15:0] _roundMask_T_16 = _GEN_0 & 16'hf0f; // @[Bitwise.scala 103:31]
  wire [15:0] _roundMask_T_18 = {_roundMask_T_11[11:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [15:0] _roundMask_T_20 = _roundMask_T_18 & 16'hf0f0; // @[Bitwise.scala 103:75]
  wire [15:0] _roundMask_T_21 = _roundMask_T_16 | _roundMask_T_20; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_1 = {{2'd0}, _roundMask_T_21[15:2]}; // @[Bitwise.scala 103:31]
  wire [15:0] _roundMask_T_26 = _GEN_1 & 16'h3333; // @[Bitwise.scala 103:31]
  wire [15:0] _roundMask_T_28 = {_roundMask_T_21[13:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [15:0] _roundMask_T_30 = _roundMask_T_28 & 16'hcccc; // @[Bitwise.scala 103:75]
  wire [15:0] _roundMask_T_31 = _roundMask_T_26 | _roundMask_T_30; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_2 = {{1'd0}, _roundMask_T_31[15:1]}; // @[Bitwise.scala 103:31]
  wire [15:0] _roundMask_T_36 = _GEN_2 & 16'h5555; // @[Bitwise.scala 103:31]
  wire [15:0] _roundMask_T_38 = {_roundMask_T_31[14:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [15:0] _roundMask_T_40 = _roundMask_T_38 & 16'haaaa; // @[Bitwise.scala 103:75]
  wire [15:0] roundMask_right = _roundMask_T_36 | _roundMask_T_40; // @[Bitwise.scala 103:39]
  wire  roundMask_right_1 = roundMask_shift[58]; // @[Bitwise.scala 109:18]
  wire  roundMask_left = roundMask_shift[59]; // @[Bitwise.scala 109:44]
  wire  roundMask_right_3 = roundMask_shift[60]; // @[Bitwise.scala 109:18]
  wire  roundMask_left_1 = roundMask_shift[61]; // @[Bitwise.scala 109:44]
  wire  roundMask_right_5 = roundMask_shift[62]; // @[Bitwise.scala 109:18]
  wire  roundMask_left_3 = roundMask_shift[63]; // @[Bitwise.scala 109:44]
  wire [21:0] _roundMask_T_46 = {roundMask_right,roundMask_right_1,roundMask_left,roundMask_right_3,roundMask_left_1,
    roundMask_right_5,roundMask_left_3}; // @[Cat.scala 29:58]
  wire [21:0] _roundMask_T_47 = ~_roundMask_T_46; // @[primitives.scala 74:36]
  wire [21:0] _roundMask_T_48 = roundMask_msb_2 ? 22'h0 : _roundMask_T_47; // @[primitives.scala 74:21]
  wire [21:0] roundMask_right_6 = ~_roundMask_T_48; // @[primitives.scala 74:17]
  wire [24:0] _roundMask_T_49 = {roundMask_right_6,3'h7}; // @[Cat.scala 29:58]
  wire  roundMask_right_7 = roundMask_shift[0]; // @[Bitwise.scala 109:18]
  wire  roundMask_left_6 = roundMask_shift[1]; // @[Bitwise.scala 109:44]
  wire  roundMask_left_7 = roundMask_shift[2]; // @[Bitwise.scala 109:44]
  wire [2:0] _roundMask_T_52 = {roundMask_right_7,roundMask_left_6,roundMask_left_7}; // @[Cat.scala 29:58]
  wire [2:0] _roundMask_T_53 = roundMask_msb_2 ? _roundMask_T_52 : 3'h0; // @[primitives.scala 61:24]
  wire [24:0] _roundMask_T_54 = roundMask_msb_1 ? _roundMask_T_49 : {{22'd0}, _roundMask_T_53}; // @[primitives.scala 66:24]
  wire [24:0] roundMask_right_9 = roundMask_msb ? _roundMask_T_54 : 25'h0; // @[primitives.scala 61:24]
  wire [26:0] roundMask = {roundMask_right_9,2'h3}; // @[Cat.scala 29:58]
  wire [25:0] shiftedRoundMask_left = roundMask[26:1]; // @[RoundAnyRawFNToRecFN.scala 160:57]
  wire [26:0] shiftedRoundMask = {1'h0,shiftedRoundMask_left}; // @[Cat.scala 29:58]
  wire [26:0] _roundPosMask_T = ~shiftedRoundMask; // @[RoundAnyRawFNToRecFN.scala 161:28]
  wire [26:0] roundPosMask = _roundPosMask_T & roundMask; // @[RoundAnyRawFNToRecFN.scala 161:46]
  wire [26:0] _roundPosBit_T = adjustedSig & roundPosMask; // @[RoundAnyRawFNToRecFN.scala 162:40]
  wire  roundPosBit = |_roundPosBit_T; // @[RoundAnyRawFNToRecFN.scala 162:56]
  wire [26:0] _anyRoundExtra_T = adjustedSig & shiftedRoundMask; // @[RoundAnyRawFNToRecFN.scala 163:42]
  wire  anyRoundExtra = |_anyRoundExtra_T; // @[RoundAnyRawFNToRecFN.scala 163:62]
  wire  anyRound = roundPosBit | anyRoundExtra; // @[RoundAnyRawFNToRecFN.scala 164:36]
  wire  _roundIncr_T = roundingMode_near_even | roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 167:38]
  wire  _roundIncr_T_1 = (roundingMode_near_even | roundingMode_near_maxMag) & roundPosBit; // @[RoundAnyRawFNToRecFN.scala 167:67]
  wire  _roundIncr_T_2 = roundMagUp & anyRound; // @[RoundAnyRawFNToRecFN.scala 169:29]
  wire  roundIncr = _roundIncr_T_1 | _roundIncr_T_2; // @[RoundAnyRawFNToRecFN.scala 168:31]
  wire [26:0] _roundedSig_T = adjustedSig | roundMask; // @[RoundAnyRawFNToRecFN.scala 172:32]
  wire [25:0] _roundedSig_T_2 = (_roundedSig_T[26:2]) + 25'h1; // @[RoundAnyRawFNToRecFN.scala 172:49]
  wire  _roundedSig_T_4 = ~anyRoundExtra; // @[RoundAnyRawFNToRecFN.scala 174:30]
  wire  _roundedSig_T_5 = (roundingMode_near_even & roundPosBit) & _roundedSig_T_4; // @[RoundAnyRawFNToRecFN.scala 173:64]
  wire [25:0] _roundedSig_T_7 = _roundedSig_T_5 ? shiftedRoundMask_left : 26'h0; // @[RoundAnyRawFNToRecFN.scala 173:25]
  wire [25:0] _roundedSig_T_8 = ~_roundedSig_T_7; // @[RoundAnyRawFNToRecFN.scala 173:21]
  wire [25:0] _roundedSig_T_9 = _roundedSig_T_2 & _roundedSig_T_8; // @[RoundAnyRawFNToRecFN.scala 172:61]
  wire [26:0] _roundedSig_T_10 = ~roundMask; // @[RoundAnyRawFNToRecFN.scala 178:32]
  wire [26:0] _roundedSig_T_11 = adjustedSig & _roundedSig_T_10; // @[RoundAnyRawFNToRecFN.scala 178:30]
  wire  _roundedSig_T_13 = roundingMode_odd & anyRound; // @[RoundAnyRawFNToRecFN.scala 179:42]
  wire [25:0] _roundedSig_T_15 = _roundedSig_T_13 ? roundPosMask[26:1] : 26'h0; // @[RoundAnyRawFNToRecFN.scala 179:24]
  wire [25:0] _GEN_3 = {{1'd0}, _roundedSig_T_11[26:2]}; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [25:0] _roundedSig_T_16 = _GEN_3 | _roundedSig_T_15; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [25:0] roundedSig = roundIncr ? _roundedSig_T_9 : _roundedSig_T_16; // @[RoundAnyRawFNToRecFN.scala 171:16]
  wire [2:0] _sRoundedExp_T_1 = {1'b0,$signed(roundedSig[25:24])}; // @[RoundAnyRawFNToRecFN.scala 183:69]
  wire [13:0] _GEN_4 = {{11{_sRoundedExp_T_1[2]}},_sRoundedExp_T_1}; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [14:0] sRoundedExp = $signed(sAdjustedExp) + $signed(_GEN_4); // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [8:0] common_expOut = sRoundedExp[8:0]; // @[RoundAnyRawFNToRecFN.scala 185:37]
  wire [22:0] common_fractOut = roundedSig[22:0]; // @[RoundAnyRawFNToRecFN.scala 189:27]
  wire [7:0] _common_overflow_T = sRoundedExp[14:7]; // @[RoundAnyRawFNToRecFN.scala 194:30]
  wire  common_overflow = $signed(_common_overflow_T) >= 8'sh3; // @[RoundAnyRawFNToRecFN.scala 194:50]
  wire  common_totalUnderflow = $signed(sRoundedExp) < 15'sh6b; // @[RoundAnyRawFNToRecFN.scala 198:31]
  wire  unboundedRange_roundPosBit = adjustedSig[1]; // @[RoundAnyRawFNToRecFN.scala 201:61]
  wire  unboundedRange_anyRound = |(adjustedSig[1:0]); // @[RoundAnyRawFNToRecFN.scala 203:70]
  wire  _unboundedRange_roundIncr_T_1 = _roundIncr_T & unboundedRange_roundPosBit; // @[RoundAnyRawFNToRecFN.scala 205:67]
  wire  _unboundedRange_roundIncr_T_2 = roundMagUp & unboundedRange_anyRound; // @[RoundAnyRawFNToRecFN.scala 207:29]
  wire  unboundedRange_roundIncr = _unboundedRange_roundIncr_T_1 | _unboundedRange_roundIncr_T_2; // @[RoundAnyRawFNToRecFN.scala 206:46]
  wire  roundCarry = roundedSig[24]; // @[RoundAnyRawFNToRecFN.scala 211:27]
  wire [5:0] _common_underflow_T = sAdjustedExp[13:8]; // @[RoundAnyRawFNToRecFN.scala 218:48]
  wire  _common_underflow_T_6 = (anyRound & ($signed(_common_underflow_T) <= 6'sh0)) & (roundMask[2]); // @[RoundAnyRawFNToRecFN.scala 218:74]
  wire  _common_underflow_T_11 = ~(roundMask[3]); // @[RoundAnyRawFNToRecFN.scala 221:34]
  wire  _common_underflow_T_13 = _common_underflow_T_11 & roundCarry; // @[RoundAnyRawFNToRecFN.scala 224:38]
  wire  _common_underflow_T_15 = (_common_underflow_T_13 & roundPosBit) & unboundedRange_roundIncr; // @[RoundAnyRawFNToRecFN.scala 225:60]
  wire  _common_underflow_T_16 = ~_common_underflow_T_15; // @[RoundAnyRawFNToRecFN.scala 220:27]
  wire  _common_underflow_T_17 = _common_underflow_T_6 & _common_underflow_T_16; // @[RoundAnyRawFNToRecFN.scala 219:76]
  wire  common_underflow = common_totalUnderflow | _common_underflow_T_17; // @[RoundAnyRawFNToRecFN.scala 215:40]
  wire  common_inexact = common_totalUnderflow | anyRound; // @[RoundAnyRawFNToRecFN.scala 228:49]
  wire  isNaNOut = io_invalidExc | io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 233:34]
  wire  commonCase = ((~isNaNOut) & (~io_in_isInf)) & (~io_in_isZero); // @[RoundAnyRawFNToRecFN.scala 235:61]
  wire  overflow = commonCase & common_overflow; // @[RoundAnyRawFNToRecFN.scala 236:32]
  wire  underflow = commonCase & common_underflow; // @[RoundAnyRawFNToRecFN.scala 237:32]
  wire  inexact = overflow | (commonCase & common_inexact); // @[RoundAnyRawFNToRecFN.scala 238:28]
  wire  overflow_roundMagUp = _roundIncr_T | roundMagUp; // @[RoundAnyRawFNToRecFN.scala 241:60]
  wire  pegMinNonzeroMagOut = (commonCase & common_totalUnderflow) & (roundMagUp | roundingMode_odd); // @[RoundAnyRawFNToRecFN.scala 243:45]
  wire  pegMaxFiniteMagOut = overflow & (~overflow_roundMagUp); // @[RoundAnyRawFNToRecFN.scala 244:39]
  wire  notNaN_isInfOut = io_in_isInf | (overflow & overflow_roundMagUp); // @[RoundAnyRawFNToRecFN.scala 246:32]
  wire  signOut = isNaNOut ? 1'h0 : io_in_sign; // @[RoundAnyRawFNToRecFN.scala 248:22]
  wire  _expOut_T = io_in_isZero | common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 251:32]
  wire [8:0] _expOut_T_1 = _expOut_T ? 9'h1c0 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 251:18]
  wire [8:0] _expOut_T_2 = ~_expOut_T_1; // @[RoundAnyRawFNToRecFN.scala 251:14]
  wire [8:0] _expOut_T_3 = common_expOut & _expOut_T_2; // @[RoundAnyRawFNToRecFN.scala 250:24]
  wire [8:0] _expOut_T_5 = pegMinNonzeroMagOut ? 9'h194 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 255:18]
  wire [8:0] _expOut_T_6 = ~_expOut_T_5; // @[RoundAnyRawFNToRecFN.scala 255:14]
  wire [8:0] _expOut_T_7 = _expOut_T_3 & _expOut_T_6; // @[RoundAnyRawFNToRecFN.scala 254:17]
  wire [8:0] _expOut_T_8 = pegMaxFiniteMagOut ? 9'h80 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 259:18]
  wire [8:0] _expOut_T_9 = ~_expOut_T_8; // @[RoundAnyRawFNToRecFN.scala 259:14]
  wire [8:0] _expOut_T_10 = _expOut_T_7 & _expOut_T_9; // @[RoundAnyRawFNToRecFN.scala 258:17]
  wire [8:0] _expOut_T_11 = notNaN_isInfOut ? 9'h40 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 263:18]
  wire [8:0] _expOut_T_12 = ~_expOut_T_11; // @[RoundAnyRawFNToRecFN.scala 263:14]
  wire [8:0] _expOut_T_13 = _expOut_T_10 & _expOut_T_12; // @[RoundAnyRawFNToRecFN.scala 262:17]
  wire [8:0] _expOut_T_14 = pegMinNonzeroMagOut ? 9'h6b : 9'h0; // @[RoundAnyRawFNToRecFN.scala 267:16]
  wire [8:0] _expOut_T_15 = _expOut_T_13 | _expOut_T_14; // @[RoundAnyRawFNToRecFN.scala 266:18]
  wire [8:0] _expOut_T_16 = pegMaxFiniteMagOut ? 9'h17f : 9'h0; // @[RoundAnyRawFNToRecFN.scala 271:16]
  wire [8:0] _expOut_T_17 = _expOut_T_15 | _expOut_T_16; // @[RoundAnyRawFNToRecFN.scala 270:15]
  wire [8:0] _expOut_T_18 = notNaN_isInfOut ? 9'h180 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 275:16]
  wire [8:0] _expOut_T_19 = _expOut_T_17 | _expOut_T_18; // @[RoundAnyRawFNToRecFN.scala 274:15]
  wire [8:0] _expOut_T_20 = isNaNOut ? 9'h1c0 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 276:16]
  wire [8:0] expOut = _expOut_T_19 | _expOut_T_20; // @[RoundAnyRawFNToRecFN.scala 275:77]
  wire  _fractOut_T_1 = (isNaNOut | io_in_isZero) | common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 278:38]
  wire [22:0] _fractOut_T_2 = isNaNOut ? 23'h400000 : 23'h0; // @[RoundAnyRawFNToRecFN.scala 279:16]
  wire [22:0] _fractOut_T_3 = _fractOut_T_1 ? _fractOut_T_2 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  wire [22:0] _fractOut_T_5 = pegMaxFiniteMagOut ? 23'h7fffff : 23'h0; // @[Bitwise.scala 72:12]
  wire [22:0] fractOut = _fractOut_T_3 | _fractOut_T_5; // @[RoundAnyRawFNToRecFN.scala 281:11]
  wire [9:0] io_out_right = {signOut,expOut}; // @[Cat.scala 29:58]
  wire [1:0] io_exceptionFlags_left = {underflow,inexact}; // @[Cat.scala 29:58]
  wire [2:0] io_exceptionFlags_right = {io_invalidExc,1'h0,overflow}; // @[Cat.scala 29:58]
  assign io_out = {io_out_right,fractOut}; // @[Cat.scala 29:58]
  assign io_exceptionFlags = {io_exceptionFlags_right,io_exceptionFlags_left}; // @[Cat.scala 29:58]
endmodule
