module DCache(
  input         gated_clock,
  input         reset,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [2:0]  auto_out_a_bits_param,
  output [3:0]  auto_out_a_bits_size,
  output        auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input  [1:0]  auto_out_b_bits_param,
  input  [3:0]  auto_out_b_bits_size,
  input         auto_out_b_bits_source,
  input  [31:0] auto_out_b_bits_address,
  input         auto_out_c_ready,
  output        auto_out_c_valid,
  output [2:0]  auto_out_c_bits_opcode,
  output [2:0]  auto_out_c_bits_param,
  output [3:0]  auto_out_c_bits_size,
  output        auto_out_c_bits_source,
  output [31:0] auto_out_c_bits_address,
  output [63:0] auto_out_c_bits_data,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [1:0]  auto_out_d_bits_param,
  input  [3:0]  auto_out_d_bits_size,
  input         auto_out_d_bits_source,
  input  [1:0]  auto_out_d_bits_sink,
  input         auto_out_d_bits_denied,
  input  [63:0] auto_out_d_bits_data,
  input         auto_out_e_ready,
  output        auto_out_e_valid,
  output [1:0]  auto_out_e_bits_sink,
  output        io_cpu_req_ready,
  input         io_cpu_req_valid,
  input  [39:0] io_cpu_req_bits_addr,
  input  [6:0]  io_cpu_req_bits_tag,
  input  [4:0]  io_cpu_req_bits_cmd,
  input  [1:0]  io_cpu_req_bits_size,
  input         io_cpu_req_bits_signed,
  input  [1:0]  io_cpu_req_bits_dprv,
  input         io_cpu_req_bits_phys,
  input         io_cpu_s1_kill,
  input  [63:0] io_cpu_s1_data_data,
  input  [7:0]  io_cpu_s1_data_mask,
  output        io_cpu_s2_nack,
  output        io_cpu_resp_valid,
  output [39:0] io_cpu_resp_bits_addr,
  output [6:0]  io_cpu_resp_bits_tag,
  output [4:0]  io_cpu_resp_bits_cmd,
  output [1:0]  io_cpu_resp_bits_size,
  output        io_cpu_resp_bits_signed,
  output [1:0]  io_cpu_resp_bits_dprv,
  output [63:0] io_cpu_resp_bits_data,
  output [7:0]  io_cpu_resp_bits_mask,
  output        io_cpu_resp_bits_replay,
  output        io_cpu_resp_bits_has_data,
  output [63:0] io_cpu_resp_bits_data_word_bypass,
  output [63:0] io_cpu_resp_bits_data_raw,
  output [63:0] io_cpu_resp_bits_store_data,
  output        io_cpu_replay_next,
  output        io_cpu_s2_xcpt_ma_ld,
  output        io_cpu_s2_xcpt_ma_st,
  output        io_cpu_s2_xcpt_pf_ld,
  output        io_cpu_s2_xcpt_pf_st,
  output        io_cpu_s2_xcpt_ae_ld,
  output        io_cpu_s2_xcpt_ae_st,
  output        io_cpu_ordered,
  output        io_cpu_perf_release,
  output        io_cpu_perf_grant,
  input         io_ptw_req_ready,
  output        io_ptw_req_valid,
  output [26:0] io_ptw_req_bits_bits_addr,
  input         io_ptw_resp_valid,
  input         io_ptw_resp_bits_ae,
  input  [53:0] io_ptw_resp_bits_pte_ppn,
  input         io_ptw_resp_bits_pte_d,
  input         io_ptw_resp_bits_pte_a,
  input         io_ptw_resp_bits_pte_g,
  input         io_ptw_resp_bits_pte_u,
  input         io_ptw_resp_bits_pte_x,
  input         io_ptw_resp_bits_pte_w,
  input         io_ptw_resp_bits_pte_r,
  input         io_ptw_resp_bits_pte_v,
  input  [1:0]  io_ptw_resp_bits_level,
  input         io_ptw_resp_bits_homogeneous,
  input  [3:0]  io_ptw_ptbr_mode,
  input         io_ptw_status_debug,
  input  [1:0]  io_ptw_status_dprv,
  input         io_ptw_status_mxr,
  input         io_ptw_status_sum,
  input         io_ptw_pmp_0_cfg_l,
  input  [1:0]  io_ptw_pmp_0_cfg_a,
  input         io_ptw_pmp_0_cfg_x,
  input         io_ptw_pmp_0_cfg_w,
  input         io_ptw_pmp_0_cfg_r,
  input  [29:0] io_ptw_pmp_0_addr,
  input  [31:0] io_ptw_pmp_0_mask,
  input         io_ptw_pmp_1_cfg_l,
  input  [1:0]  io_ptw_pmp_1_cfg_a,
  input         io_ptw_pmp_1_cfg_x,
  input         io_ptw_pmp_1_cfg_w,
  input         io_ptw_pmp_1_cfg_r,
  input  [29:0] io_ptw_pmp_1_addr,
  input  [31:0] io_ptw_pmp_1_mask,
  input         io_ptw_pmp_2_cfg_l,
  input  [1:0]  io_ptw_pmp_2_cfg_a,
  input         io_ptw_pmp_2_cfg_x,
  input         io_ptw_pmp_2_cfg_w,
  input         io_ptw_pmp_2_cfg_r,
  input  [29:0] io_ptw_pmp_2_addr,
  input  [31:0] io_ptw_pmp_2_mask,
  input         io_ptw_pmp_3_cfg_l,
  input  [1:0]  io_ptw_pmp_3_cfg_a,
  input         io_ptw_pmp_3_cfg_x,
  input         io_ptw_pmp_3_cfg_w,
  input         io_ptw_pmp_3_cfg_r,
  input  [29:0] io_ptw_pmp_3_addr,
  input  [31:0] io_ptw_pmp_3_mask,
  input         io_ptw_pmp_4_cfg_l,
  input  [1:0]  io_ptw_pmp_4_cfg_a,
  input         io_ptw_pmp_4_cfg_x,
  input         io_ptw_pmp_4_cfg_w,
  input         io_ptw_pmp_4_cfg_r,
  input  [29:0] io_ptw_pmp_4_addr,
  input  [31:0] io_ptw_pmp_4_mask,
  input         io_ptw_pmp_5_cfg_l,
  input  [1:0]  io_ptw_pmp_5_cfg_a,
  input         io_ptw_pmp_5_cfg_x,
  input         io_ptw_pmp_5_cfg_w,
  input         io_ptw_pmp_5_cfg_r,
  input  [29:0] io_ptw_pmp_5_addr,
  input  [31:0] io_ptw_pmp_5_mask,
  input         io_ptw_pmp_6_cfg_l,
  input  [1:0]  io_ptw_pmp_6_cfg_a,
  input         io_ptw_pmp_6_cfg_x,
  input         io_ptw_pmp_6_cfg_w,
  input         io_ptw_pmp_6_cfg_r,
  input  [29:0] io_ptw_pmp_6_addr,
  input  [31:0] io_ptw_pmp_6_mask,
  input         io_ptw_pmp_7_cfg_l,
  input  [1:0]  io_ptw_pmp_7_cfg_a,
  input         io_ptw_pmp_7_cfg_x,
  input         io_ptw_pmp_7_cfg_w,
  input         io_ptw_pmp_7_cfg_r,
  input  [29:0] io_ptw_pmp_7_addr,
  input  [31:0] io_ptw_pmp_7_mask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [63:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [63:0] _RAND_120;
  reg [63:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [63:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [63:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [63:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [63:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [63:0] _RAND_158;
  reg [63:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [63:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [63:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [63:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
`endif // RANDOMIZE_REG_INIT
  wire  tlb_clock;
  wire  tlb_reset;
  wire  tlb_io_req_ready;
  wire  tlb_io_req_valid;
  wire [39:0] tlb_io_req_bits_vaddr;
  wire  tlb_io_req_bits_passthrough;
  wire [1:0] tlb_io_req_bits_size;
  wire [4:0] tlb_io_req_bits_cmd;
  wire  tlb_io_resp_miss;
  wire [31:0] tlb_io_resp_paddr;
  wire  tlb_io_resp_pf_ld;
  wire  tlb_io_resp_pf_st;
  wire  tlb_io_resp_ae_ld;
  wire  tlb_io_resp_ae_st;
  wire  tlb_io_resp_ma_ld;
  wire  tlb_io_resp_ma_st;
  wire  tlb_io_resp_cacheable;
  wire  tlb_io_sfence_valid;
  wire  tlb_io_sfence_bits_rs1;
  wire  tlb_io_sfence_bits_rs2;
  wire [38:0] tlb_io_sfence_bits_addr;
  wire  tlb_io_ptw_req_ready;
  wire  tlb_io_ptw_req_valid;
  wire [26:0] tlb_io_ptw_req_bits_bits_addr;
  wire  tlb_io_ptw_resp_valid;
  wire  tlb_io_ptw_resp_bits_ae;
  wire [53:0] tlb_io_ptw_resp_bits_pte_ppn;
  wire  tlb_io_ptw_resp_bits_pte_d;
  wire  tlb_io_ptw_resp_bits_pte_a;
  wire  tlb_io_ptw_resp_bits_pte_g;
  wire  tlb_io_ptw_resp_bits_pte_u;
  wire  tlb_io_ptw_resp_bits_pte_x;
  wire  tlb_io_ptw_resp_bits_pte_w;
  wire  tlb_io_ptw_resp_bits_pte_r;
  wire  tlb_io_ptw_resp_bits_pte_v;
  wire [1:0] tlb_io_ptw_resp_bits_level;
  wire  tlb_io_ptw_resp_bits_homogeneous;
  wire [3:0] tlb_io_ptw_ptbr_mode;
  wire  tlb_io_ptw_status_debug;
  wire [1:0] tlb_io_ptw_status_dprv;
  wire  tlb_io_ptw_status_mxr;
  wire  tlb_io_ptw_status_sum;
  wire  tlb_io_ptw_pmp_0_cfg_l;
  wire [1:0] tlb_io_ptw_pmp_0_cfg_a;
  wire  tlb_io_ptw_pmp_0_cfg_x;
  wire  tlb_io_ptw_pmp_0_cfg_w;
  wire  tlb_io_ptw_pmp_0_cfg_r;
  wire [29:0] tlb_io_ptw_pmp_0_addr;
  wire [31:0] tlb_io_ptw_pmp_0_mask;
  wire  tlb_io_ptw_pmp_1_cfg_l;
  wire [1:0] tlb_io_ptw_pmp_1_cfg_a;
  wire  tlb_io_ptw_pmp_1_cfg_x;
  wire  tlb_io_ptw_pmp_1_cfg_w;
  wire  tlb_io_ptw_pmp_1_cfg_r;
  wire [29:0] tlb_io_ptw_pmp_1_addr;
  wire [31:0] tlb_io_ptw_pmp_1_mask;
  wire  tlb_io_ptw_pmp_2_cfg_l;
  wire [1:0] tlb_io_ptw_pmp_2_cfg_a;
  wire  tlb_io_ptw_pmp_2_cfg_x;
  wire  tlb_io_ptw_pmp_2_cfg_w;
  wire  tlb_io_ptw_pmp_2_cfg_r;
  wire [29:0] tlb_io_ptw_pmp_2_addr;
  wire [31:0] tlb_io_ptw_pmp_2_mask;
  wire  tlb_io_ptw_pmp_3_cfg_l;
  wire [1:0] tlb_io_ptw_pmp_3_cfg_a;
  wire  tlb_io_ptw_pmp_3_cfg_x;
  wire  tlb_io_ptw_pmp_3_cfg_w;
  wire  tlb_io_ptw_pmp_3_cfg_r;
  wire [29:0] tlb_io_ptw_pmp_3_addr;
  wire [31:0] tlb_io_ptw_pmp_3_mask;
  wire  tlb_io_ptw_pmp_4_cfg_l;
  wire [1:0] tlb_io_ptw_pmp_4_cfg_a;
  wire  tlb_io_ptw_pmp_4_cfg_x;
  wire  tlb_io_ptw_pmp_4_cfg_w;
  wire  tlb_io_ptw_pmp_4_cfg_r;
  wire [29:0] tlb_io_ptw_pmp_4_addr;
  wire [31:0] tlb_io_ptw_pmp_4_mask;
  wire  tlb_io_ptw_pmp_5_cfg_l;
  wire [1:0] tlb_io_ptw_pmp_5_cfg_a;
  wire  tlb_io_ptw_pmp_5_cfg_x;
  wire  tlb_io_ptw_pmp_5_cfg_w;
  wire  tlb_io_ptw_pmp_5_cfg_r;
  wire [29:0] tlb_io_ptw_pmp_5_addr;
  wire [31:0] tlb_io_ptw_pmp_5_mask;
  wire  tlb_io_ptw_pmp_6_cfg_l;
  wire [1:0] tlb_io_ptw_pmp_6_cfg_a;
  wire  tlb_io_ptw_pmp_6_cfg_x;
  wire  tlb_io_ptw_pmp_6_cfg_w;
  wire  tlb_io_ptw_pmp_6_cfg_r;
  wire [29:0] tlb_io_ptw_pmp_6_addr;
  wire [31:0] tlb_io_ptw_pmp_6_mask;
  wire  tlb_io_ptw_pmp_7_cfg_l;
  wire [1:0] tlb_io_ptw_pmp_7_cfg_a;
  wire  tlb_io_ptw_pmp_7_cfg_x;
  wire  tlb_io_ptw_pmp_7_cfg_w;
  wire  tlb_io_ptw_pmp_7_cfg_r;
  wire [29:0] tlb_io_ptw_pmp_7_addr;
  wire [31:0] tlb_io_ptw_pmp_7_mask;
  wire [19:0] tlb_mpu_ppn_data_barrier_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_mpu_ppn_data_barrier_io_x_u; // @[package.scala 236:25]
  wire  tlb_mpu_ppn_data_barrier_io_x_ae; // @[package.scala 236:25]
  wire  tlb_mpu_ppn_data_barrier_io_x_sw; // @[package.scala 236:25]
  wire  tlb_mpu_ppn_data_barrier_io_x_sx; // @[package.scala 236:25]
  wire  tlb_mpu_ppn_data_barrier_io_x_sr; // @[package.scala 236:25]
  wire  tlb_mpu_ppn_data_barrier_io_x_pw; // @[package.scala 236:25]
  wire  tlb_mpu_ppn_data_barrier_io_x_px; // @[package.scala 236:25]
  wire  tlb_mpu_ppn_data_barrier_io_x_pr; // @[package.scala 236:25]
  wire  tlb_mpu_ppn_data_barrier_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_mpu_ppn_data_barrier_io_x_pal; // @[package.scala 236:25]
  wire  tlb_mpu_ppn_data_barrier_io_x_paa; // @[package.scala 236:25]
  wire  tlb_mpu_ppn_data_barrier_io_x_eff; // @[package.scala 236:25]
  wire  tlb_mpu_ppn_data_barrier_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_mpu_ppn_data_barrier_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_mpu_ppn_data_barrier_io_y_u; // @[package.scala 236:25]
  wire  tlb_mpu_ppn_data_barrier_io_y_ae; // @[package.scala 236:25]
  wire  tlb_mpu_ppn_data_barrier_io_y_sw; // @[package.scala 236:25]
  wire  tlb_mpu_ppn_data_barrier_io_y_sx; // @[package.scala 236:25]
  wire  tlb_mpu_ppn_data_barrier_io_y_sr; // @[package.scala 236:25]
  wire  tlb_mpu_ppn_data_barrier_io_y_pw; // @[package.scala 236:25]
  wire  tlb_mpu_ppn_data_barrier_io_y_px; // @[package.scala 236:25]
  wire  tlb_mpu_ppn_data_barrier_io_y_pr; // @[package.scala 236:25]
  wire  tlb_mpu_ppn_data_barrier_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_mpu_ppn_data_barrier_io_y_pal; // @[package.scala 236:25]
  wire  tlb_mpu_ppn_data_barrier_io_y_paa; // @[package.scala 236:25]
  wire  tlb_mpu_ppn_data_barrier_io_y_eff; // @[package.scala 236:25]
  wire  tlb_mpu_ppn_data_barrier_io_y_c; // @[package.scala 236:25]
  wire [1:0] tlb_pmp_io_prv; // @[TLB.scala 190:19]
  wire  tlb_pmp_io_pmp_0_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] tlb_pmp_io_pmp_0_cfg_a; // @[TLB.scala 190:19]
  wire  tlb_pmp_io_pmp_0_cfg_x; // @[TLB.scala 190:19]
  wire  tlb_pmp_io_pmp_0_cfg_w; // @[TLB.scala 190:19]
  wire  tlb_pmp_io_pmp_0_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] tlb_pmp_io_pmp_0_addr; // @[TLB.scala 190:19]
  wire [31:0] tlb_pmp_io_pmp_0_mask; // @[TLB.scala 190:19]
  wire  tlb_pmp_io_pmp_1_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] tlb_pmp_io_pmp_1_cfg_a; // @[TLB.scala 190:19]
  wire  tlb_pmp_io_pmp_1_cfg_x; // @[TLB.scala 190:19]
  wire  tlb_pmp_io_pmp_1_cfg_w; // @[TLB.scala 190:19]
  wire  tlb_pmp_io_pmp_1_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] tlb_pmp_io_pmp_1_addr; // @[TLB.scala 190:19]
  wire [31:0] tlb_pmp_io_pmp_1_mask; // @[TLB.scala 190:19]
  wire  tlb_pmp_io_pmp_2_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] tlb_pmp_io_pmp_2_cfg_a; // @[TLB.scala 190:19]
  wire  tlb_pmp_io_pmp_2_cfg_x; // @[TLB.scala 190:19]
  wire  tlb_pmp_io_pmp_2_cfg_w; // @[TLB.scala 190:19]
  wire  tlb_pmp_io_pmp_2_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] tlb_pmp_io_pmp_2_addr; // @[TLB.scala 190:19]
  wire [31:0] tlb_pmp_io_pmp_2_mask; // @[TLB.scala 190:19]
  wire  tlb_pmp_io_pmp_3_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] tlb_pmp_io_pmp_3_cfg_a; // @[TLB.scala 190:19]
  wire  tlb_pmp_io_pmp_3_cfg_x; // @[TLB.scala 190:19]
  wire  tlb_pmp_io_pmp_3_cfg_w; // @[TLB.scala 190:19]
  wire  tlb_pmp_io_pmp_3_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] tlb_pmp_io_pmp_3_addr; // @[TLB.scala 190:19]
  wire [31:0] tlb_pmp_io_pmp_3_mask; // @[TLB.scala 190:19]
  wire  tlb_pmp_io_pmp_4_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] tlb_pmp_io_pmp_4_cfg_a; // @[TLB.scala 190:19]
  wire  tlb_pmp_io_pmp_4_cfg_x; // @[TLB.scala 190:19]
  wire  tlb_pmp_io_pmp_4_cfg_w; // @[TLB.scala 190:19]
  wire  tlb_pmp_io_pmp_4_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] tlb_pmp_io_pmp_4_addr; // @[TLB.scala 190:19]
  wire [31:0] tlb_pmp_io_pmp_4_mask; // @[TLB.scala 190:19]
  wire  tlb_pmp_io_pmp_5_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] tlb_pmp_io_pmp_5_cfg_a; // @[TLB.scala 190:19]
  wire  tlb_pmp_io_pmp_5_cfg_x; // @[TLB.scala 190:19]
  wire  tlb_pmp_io_pmp_5_cfg_w; // @[TLB.scala 190:19]
  wire  tlb_pmp_io_pmp_5_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] tlb_pmp_io_pmp_5_addr; // @[TLB.scala 190:19]
  wire [31:0] tlb_pmp_io_pmp_5_mask; // @[TLB.scala 190:19]
  wire  tlb_pmp_io_pmp_6_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] tlb_pmp_io_pmp_6_cfg_a; // @[TLB.scala 190:19]
  wire  tlb_pmp_io_pmp_6_cfg_x; // @[TLB.scala 190:19]
  wire  tlb_pmp_io_pmp_6_cfg_w; // @[TLB.scala 190:19]
  wire  tlb_pmp_io_pmp_6_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] tlb_pmp_io_pmp_6_addr; // @[TLB.scala 190:19]
  wire [31:0] tlb_pmp_io_pmp_6_mask; // @[TLB.scala 190:19]
  wire  tlb_pmp_io_pmp_7_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] tlb_pmp_io_pmp_7_cfg_a; // @[TLB.scala 190:19]
  wire  tlb_pmp_io_pmp_7_cfg_x; // @[TLB.scala 190:19]
  wire  tlb_pmp_io_pmp_7_cfg_w; // @[TLB.scala 190:19]
  wire  tlb_pmp_io_pmp_7_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] tlb_pmp_io_pmp_7_addr; // @[TLB.scala 190:19]
  wire [31:0] tlb_pmp_io_pmp_7_mask; // @[TLB.scala 190:19]
  wire [31:0] tlb_pmp_io_addr; // @[TLB.scala 190:19]
  wire [1:0] tlb_pmp_io_size; // @[TLB.scala 190:19]
  wire  tlb_pmp_io_r; // @[TLB.scala 190:19]
  wire  tlb_pmp_io_w; // @[TLB.scala 190:19]
  wire  tlb_pmp_io_x; // @[TLB.scala 190:19]
  wire [19:0] tlb_ppn_data_barrier_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_io_x_u; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_io_x_ae; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_io_x_sw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_io_x_sx; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_io_x_sr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_io_x_pw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_io_x_px; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_io_x_pr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_io_x_pal; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_io_x_paa; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_io_x_eff; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_ppn_data_barrier_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_io_y_u; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_io_y_ae; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_io_y_sw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_io_y_sx; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_io_y_sr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_io_y_pw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_io_y_px; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_io_y_pr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_io_y_pal; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_io_y_paa; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_io_y_eff; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_ppn_data_barrier_1_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_1_io_x_u; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_1_io_x_ae; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_1_io_x_sw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_1_io_x_sx; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_1_io_x_sr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_1_io_x_pw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_1_io_x_px; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_1_io_x_pr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_1_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_1_io_x_pal; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_1_io_x_paa; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_1_io_x_eff; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_1_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_ppn_data_barrier_1_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_1_io_y_u; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_1_io_y_ae; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_1_io_y_sw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_1_io_y_sx; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_1_io_y_sr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_1_io_y_pw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_1_io_y_px; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_1_io_y_pr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_1_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_1_io_y_pal; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_1_io_y_paa; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_1_io_y_eff; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_1_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_ppn_data_barrier_2_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_2_io_x_u; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_2_io_x_ae; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_2_io_x_sw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_2_io_x_sx; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_2_io_x_sr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_2_io_x_pw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_2_io_x_px; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_2_io_x_pr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_2_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_2_io_x_pal; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_2_io_x_paa; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_2_io_x_eff; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_2_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_ppn_data_barrier_2_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_2_io_y_u; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_2_io_y_ae; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_2_io_y_sw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_2_io_y_sx; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_2_io_y_sr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_2_io_y_pw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_2_io_y_px; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_2_io_y_pr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_2_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_2_io_y_pal; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_2_io_y_paa; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_2_io_y_eff; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_2_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_ppn_data_barrier_3_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_3_io_x_u; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_3_io_x_ae; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_3_io_x_sw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_3_io_x_sx; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_3_io_x_sr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_3_io_x_pw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_3_io_x_px; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_3_io_x_pr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_3_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_3_io_x_pal; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_3_io_x_paa; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_3_io_x_eff; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_3_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_ppn_data_barrier_3_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_3_io_y_u; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_3_io_y_ae; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_3_io_y_sw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_3_io_y_sx; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_3_io_y_sr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_3_io_y_pw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_3_io_y_px; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_3_io_y_pr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_3_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_3_io_y_pal; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_3_io_y_paa; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_3_io_y_eff; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_3_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_ppn_data_barrier_4_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_4_io_x_u; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_4_io_x_ae; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_4_io_x_sw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_4_io_x_sx; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_4_io_x_sr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_4_io_x_pw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_4_io_x_px; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_4_io_x_pr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_4_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_4_io_x_pal; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_4_io_x_paa; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_4_io_x_eff; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_4_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_ppn_data_barrier_4_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_4_io_y_u; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_4_io_y_ae; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_4_io_y_sw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_4_io_y_sx; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_4_io_y_sr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_4_io_y_pw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_4_io_y_px; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_4_io_y_pr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_4_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_4_io_y_pal; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_4_io_y_paa; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_4_io_y_eff; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_4_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_ppn_data_barrier_5_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_5_io_x_u; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_5_io_x_ae; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_5_io_x_sw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_5_io_x_sx; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_5_io_x_sr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_5_io_x_pw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_5_io_x_px; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_5_io_x_pr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_5_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_5_io_x_pal; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_5_io_x_paa; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_5_io_x_eff; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_5_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_ppn_data_barrier_5_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_5_io_y_u; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_5_io_y_ae; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_5_io_y_sw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_5_io_y_sx; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_5_io_y_sr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_5_io_y_pw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_5_io_y_px; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_5_io_y_pr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_5_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_5_io_y_pal; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_5_io_y_paa; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_5_io_y_eff; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_5_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_ppn_data_barrier_6_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_6_io_x_u; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_6_io_x_ae; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_6_io_x_sw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_6_io_x_sx; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_6_io_x_sr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_6_io_x_pw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_6_io_x_px; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_6_io_x_pr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_6_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_6_io_x_pal; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_6_io_x_paa; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_6_io_x_eff; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_6_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_ppn_data_barrier_6_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_6_io_y_u; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_6_io_y_ae; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_6_io_y_sw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_6_io_y_sx; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_6_io_y_sr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_6_io_y_pw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_6_io_y_px; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_6_io_y_pr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_6_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_6_io_y_pal; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_6_io_y_paa; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_6_io_y_eff; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_6_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_ppn_data_barrier_7_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_7_io_x_u; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_7_io_x_ae; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_7_io_x_sw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_7_io_x_sx; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_7_io_x_sr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_7_io_x_pw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_7_io_x_px; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_7_io_x_pr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_7_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_7_io_x_pal; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_7_io_x_paa; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_7_io_x_eff; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_7_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_ppn_data_barrier_7_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_7_io_y_u; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_7_io_y_ae; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_7_io_y_sw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_7_io_y_sx; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_7_io_y_sr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_7_io_y_pw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_7_io_y_px; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_7_io_y_pr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_7_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_7_io_y_pal; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_7_io_y_paa; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_7_io_y_eff; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_7_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_ppn_data_barrier_8_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_8_io_x_u; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_8_io_x_ae; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_8_io_x_sw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_8_io_x_sx; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_8_io_x_sr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_8_io_x_pw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_8_io_x_px; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_8_io_x_pr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_8_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_8_io_x_pal; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_8_io_x_paa; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_8_io_x_eff; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_8_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_ppn_data_barrier_8_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_8_io_y_u; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_8_io_y_ae; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_8_io_y_sw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_8_io_y_sx; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_8_io_y_sr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_8_io_y_pw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_8_io_y_px; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_8_io_y_pr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_8_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_8_io_y_pal; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_8_io_y_paa; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_8_io_y_eff; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_8_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_ppn_data_barrier_9_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_9_io_x_u; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_9_io_x_ae; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_9_io_x_sw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_9_io_x_sx; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_9_io_x_sr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_9_io_x_pw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_9_io_x_px; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_9_io_x_pr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_9_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_9_io_x_pal; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_9_io_x_paa; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_9_io_x_eff; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_9_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_ppn_data_barrier_9_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_9_io_y_u; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_9_io_y_ae; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_9_io_y_sw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_9_io_y_sx; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_9_io_y_sr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_9_io_y_pw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_9_io_y_px; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_9_io_y_pr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_9_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_9_io_y_pal; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_9_io_y_paa; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_9_io_y_eff; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_9_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_ppn_data_barrier_10_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_10_io_x_u; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_10_io_x_ae; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_10_io_x_sw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_10_io_x_sx; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_10_io_x_sr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_10_io_x_pw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_10_io_x_px; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_10_io_x_pr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_10_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_10_io_x_pal; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_10_io_x_paa; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_10_io_x_eff; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_10_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_ppn_data_barrier_10_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_10_io_y_u; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_10_io_y_ae; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_10_io_y_sw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_10_io_y_sx; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_10_io_y_sr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_10_io_y_pw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_10_io_y_px; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_10_io_y_pr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_10_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_10_io_y_pal; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_10_io_y_paa; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_10_io_y_eff; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_10_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_ppn_data_barrier_11_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_11_io_x_u; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_11_io_x_ae; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_11_io_x_sw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_11_io_x_sx; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_11_io_x_sr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_11_io_x_pw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_11_io_x_px; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_11_io_x_pr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_11_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_11_io_x_pal; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_11_io_x_paa; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_11_io_x_eff; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_11_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_ppn_data_barrier_11_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_11_io_y_u; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_11_io_y_ae; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_11_io_y_sw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_11_io_y_sx; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_11_io_y_sr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_11_io_y_pw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_11_io_y_px; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_11_io_y_pr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_11_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_11_io_y_pal; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_11_io_y_paa; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_11_io_y_eff; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_11_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_ppn_data_barrier_12_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_12_io_x_u; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_12_io_x_ae; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_12_io_x_sw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_12_io_x_sx; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_12_io_x_sr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_12_io_x_pw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_12_io_x_px; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_12_io_x_pr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_12_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_12_io_x_pal; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_12_io_x_paa; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_12_io_x_eff; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_12_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_ppn_data_barrier_12_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_12_io_y_u; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_12_io_y_ae; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_12_io_y_sw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_12_io_y_sx; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_12_io_y_sr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_12_io_y_pw; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_12_io_y_px; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_12_io_y_pr; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_12_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_12_io_y_pal; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_12_io_y_paa; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_12_io_y_eff; // @[package.scala 236:25]
  wire  tlb_ppn_data_barrier_12_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_entries_barrier_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_entries_barrier_io_x_u; // @[package.scala 236:25]
  wire  tlb_entries_barrier_io_x_ae; // @[package.scala 236:25]
  wire  tlb_entries_barrier_io_x_sw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_io_x_sx; // @[package.scala 236:25]
  wire  tlb_entries_barrier_io_x_sr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_io_x_pw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_io_x_px; // @[package.scala 236:25]
  wire  tlb_entries_barrier_io_x_pr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_entries_barrier_io_x_pal; // @[package.scala 236:25]
  wire  tlb_entries_barrier_io_x_paa; // @[package.scala 236:25]
  wire  tlb_entries_barrier_io_x_eff; // @[package.scala 236:25]
  wire  tlb_entries_barrier_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_entries_barrier_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_entries_barrier_io_y_u; // @[package.scala 236:25]
  wire  tlb_entries_barrier_io_y_ae; // @[package.scala 236:25]
  wire  tlb_entries_barrier_io_y_sw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_io_y_sx; // @[package.scala 236:25]
  wire  tlb_entries_barrier_io_y_sr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_io_y_pw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_io_y_px; // @[package.scala 236:25]
  wire  tlb_entries_barrier_io_y_pr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_entries_barrier_io_y_pal; // @[package.scala 236:25]
  wire  tlb_entries_barrier_io_y_paa; // @[package.scala 236:25]
  wire  tlb_entries_barrier_io_y_eff; // @[package.scala 236:25]
  wire  tlb_entries_barrier_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_entries_barrier_1_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_entries_barrier_1_io_x_u; // @[package.scala 236:25]
  wire  tlb_entries_barrier_1_io_x_ae; // @[package.scala 236:25]
  wire  tlb_entries_barrier_1_io_x_sw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_1_io_x_sx; // @[package.scala 236:25]
  wire  tlb_entries_barrier_1_io_x_sr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_1_io_x_pw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_1_io_x_px; // @[package.scala 236:25]
  wire  tlb_entries_barrier_1_io_x_pr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_1_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_entries_barrier_1_io_x_pal; // @[package.scala 236:25]
  wire  tlb_entries_barrier_1_io_x_paa; // @[package.scala 236:25]
  wire  tlb_entries_barrier_1_io_x_eff; // @[package.scala 236:25]
  wire  tlb_entries_barrier_1_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_entries_barrier_1_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_entries_barrier_1_io_y_u; // @[package.scala 236:25]
  wire  tlb_entries_barrier_1_io_y_ae; // @[package.scala 236:25]
  wire  tlb_entries_barrier_1_io_y_sw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_1_io_y_sx; // @[package.scala 236:25]
  wire  tlb_entries_barrier_1_io_y_sr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_1_io_y_pw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_1_io_y_px; // @[package.scala 236:25]
  wire  tlb_entries_barrier_1_io_y_pr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_1_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_entries_barrier_1_io_y_pal; // @[package.scala 236:25]
  wire  tlb_entries_barrier_1_io_y_paa; // @[package.scala 236:25]
  wire  tlb_entries_barrier_1_io_y_eff; // @[package.scala 236:25]
  wire  tlb_entries_barrier_1_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_entries_barrier_2_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_entries_barrier_2_io_x_u; // @[package.scala 236:25]
  wire  tlb_entries_barrier_2_io_x_ae; // @[package.scala 236:25]
  wire  tlb_entries_barrier_2_io_x_sw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_2_io_x_sx; // @[package.scala 236:25]
  wire  tlb_entries_barrier_2_io_x_sr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_2_io_x_pw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_2_io_x_px; // @[package.scala 236:25]
  wire  tlb_entries_barrier_2_io_x_pr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_2_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_entries_barrier_2_io_x_pal; // @[package.scala 236:25]
  wire  tlb_entries_barrier_2_io_x_paa; // @[package.scala 236:25]
  wire  tlb_entries_barrier_2_io_x_eff; // @[package.scala 236:25]
  wire  tlb_entries_barrier_2_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_entries_barrier_2_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_entries_barrier_2_io_y_u; // @[package.scala 236:25]
  wire  tlb_entries_barrier_2_io_y_ae; // @[package.scala 236:25]
  wire  tlb_entries_barrier_2_io_y_sw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_2_io_y_sx; // @[package.scala 236:25]
  wire  tlb_entries_barrier_2_io_y_sr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_2_io_y_pw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_2_io_y_px; // @[package.scala 236:25]
  wire  tlb_entries_barrier_2_io_y_pr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_2_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_entries_barrier_2_io_y_pal; // @[package.scala 236:25]
  wire  tlb_entries_barrier_2_io_y_paa; // @[package.scala 236:25]
  wire  tlb_entries_barrier_2_io_y_eff; // @[package.scala 236:25]
  wire  tlb_entries_barrier_2_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_entries_barrier_3_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_entries_barrier_3_io_x_u; // @[package.scala 236:25]
  wire  tlb_entries_barrier_3_io_x_ae; // @[package.scala 236:25]
  wire  tlb_entries_barrier_3_io_x_sw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_3_io_x_sx; // @[package.scala 236:25]
  wire  tlb_entries_barrier_3_io_x_sr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_3_io_x_pw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_3_io_x_px; // @[package.scala 236:25]
  wire  tlb_entries_barrier_3_io_x_pr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_3_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_entries_barrier_3_io_x_pal; // @[package.scala 236:25]
  wire  tlb_entries_barrier_3_io_x_paa; // @[package.scala 236:25]
  wire  tlb_entries_barrier_3_io_x_eff; // @[package.scala 236:25]
  wire  tlb_entries_barrier_3_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_entries_barrier_3_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_entries_barrier_3_io_y_u; // @[package.scala 236:25]
  wire  tlb_entries_barrier_3_io_y_ae; // @[package.scala 236:25]
  wire  tlb_entries_barrier_3_io_y_sw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_3_io_y_sx; // @[package.scala 236:25]
  wire  tlb_entries_barrier_3_io_y_sr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_3_io_y_pw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_3_io_y_px; // @[package.scala 236:25]
  wire  tlb_entries_barrier_3_io_y_pr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_3_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_entries_barrier_3_io_y_pal; // @[package.scala 236:25]
  wire  tlb_entries_barrier_3_io_y_paa; // @[package.scala 236:25]
  wire  tlb_entries_barrier_3_io_y_eff; // @[package.scala 236:25]
  wire  tlb_entries_barrier_3_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_entries_barrier_4_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_entries_barrier_4_io_x_u; // @[package.scala 236:25]
  wire  tlb_entries_barrier_4_io_x_ae; // @[package.scala 236:25]
  wire  tlb_entries_barrier_4_io_x_sw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_4_io_x_sx; // @[package.scala 236:25]
  wire  tlb_entries_barrier_4_io_x_sr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_4_io_x_pw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_4_io_x_px; // @[package.scala 236:25]
  wire  tlb_entries_barrier_4_io_x_pr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_4_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_entries_barrier_4_io_x_pal; // @[package.scala 236:25]
  wire  tlb_entries_barrier_4_io_x_paa; // @[package.scala 236:25]
  wire  tlb_entries_barrier_4_io_x_eff; // @[package.scala 236:25]
  wire  tlb_entries_barrier_4_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_entries_barrier_4_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_entries_barrier_4_io_y_u; // @[package.scala 236:25]
  wire  tlb_entries_barrier_4_io_y_ae; // @[package.scala 236:25]
  wire  tlb_entries_barrier_4_io_y_sw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_4_io_y_sx; // @[package.scala 236:25]
  wire  tlb_entries_barrier_4_io_y_sr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_4_io_y_pw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_4_io_y_px; // @[package.scala 236:25]
  wire  tlb_entries_barrier_4_io_y_pr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_4_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_entries_barrier_4_io_y_pal; // @[package.scala 236:25]
  wire  tlb_entries_barrier_4_io_y_paa; // @[package.scala 236:25]
  wire  tlb_entries_barrier_4_io_y_eff; // @[package.scala 236:25]
  wire  tlb_entries_barrier_4_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_entries_barrier_5_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_entries_barrier_5_io_x_u; // @[package.scala 236:25]
  wire  tlb_entries_barrier_5_io_x_ae; // @[package.scala 236:25]
  wire  tlb_entries_barrier_5_io_x_sw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_5_io_x_sx; // @[package.scala 236:25]
  wire  tlb_entries_barrier_5_io_x_sr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_5_io_x_pw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_5_io_x_px; // @[package.scala 236:25]
  wire  tlb_entries_barrier_5_io_x_pr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_5_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_entries_barrier_5_io_x_pal; // @[package.scala 236:25]
  wire  tlb_entries_barrier_5_io_x_paa; // @[package.scala 236:25]
  wire  tlb_entries_barrier_5_io_x_eff; // @[package.scala 236:25]
  wire  tlb_entries_barrier_5_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_entries_barrier_5_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_entries_barrier_5_io_y_u; // @[package.scala 236:25]
  wire  tlb_entries_barrier_5_io_y_ae; // @[package.scala 236:25]
  wire  tlb_entries_barrier_5_io_y_sw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_5_io_y_sx; // @[package.scala 236:25]
  wire  tlb_entries_barrier_5_io_y_sr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_5_io_y_pw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_5_io_y_px; // @[package.scala 236:25]
  wire  tlb_entries_barrier_5_io_y_pr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_5_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_entries_barrier_5_io_y_pal; // @[package.scala 236:25]
  wire  tlb_entries_barrier_5_io_y_paa; // @[package.scala 236:25]
  wire  tlb_entries_barrier_5_io_y_eff; // @[package.scala 236:25]
  wire  tlb_entries_barrier_5_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_entries_barrier_6_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_entries_barrier_6_io_x_u; // @[package.scala 236:25]
  wire  tlb_entries_barrier_6_io_x_ae; // @[package.scala 236:25]
  wire  tlb_entries_barrier_6_io_x_sw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_6_io_x_sx; // @[package.scala 236:25]
  wire  tlb_entries_barrier_6_io_x_sr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_6_io_x_pw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_6_io_x_px; // @[package.scala 236:25]
  wire  tlb_entries_barrier_6_io_x_pr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_6_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_entries_barrier_6_io_x_pal; // @[package.scala 236:25]
  wire  tlb_entries_barrier_6_io_x_paa; // @[package.scala 236:25]
  wire  tlb_entries_barrier_6_io_x_eff; // @[package.scala 236:25]
  wire  tlb_entries_barrier_6_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_entries_barrier_6_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_entries_barrier_6_io_y_u; // @[package.scala 236:25]
  wire  tlb_entries_barrier_6_io_y_ae; // @[package.scala 236:25]
  wire  tlb_entries_barrier_6_io_y_sw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_6_io_y_sx; // @[package.scala 236:25]
  wire  tlb_entries_barrier_6_io_y_sr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_6_io_y_pw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_6_io_y_px; // @[package.scala 236:25]
  wire  tlb_entries_barrier_6_io_y_pr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_6_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_entries_barrier_6_io_y_pal; // @[package.scala 236:25]
  wire  tlb_entries_barrier_6_io_y_paa; // @[package.scala 236:25]
  wire  tlb_entries_barrier_6_io_y_eff; // @[package.scala 236:25]
  wire  tlb_entries_barrier_6_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_entries_barrier_7_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_entries_barrier_7_io_x_u; // @[package.scala 236:25]
  wire  tlb_entries_barrier_7_io_x_ae; // @[package.scala 236:25]
  wire  tlb_entries_barrier_7_io_x_sw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_7_io_x_sx; // @[package.scala 236:25]
  wire  tlb_entries_barrier_7_io_x_sr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_7_io_x_pw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_7_io_x_px; // @[package.scala 236:25]
  wire  tlb_entries_barrier_7_io_x_pr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_7_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_entries_barrier_7_io_x_pal; // @[package.scala 236:25]
  wire  tlb_entries_barrier_7_io_x_paa; // @[package.scala 236:25]
  wire  tlb_entries_barrier_7_io_x_eff; // @[package.scala 236:25]
  wire  tlb_entries_barrier_7_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_entries_barrier_7_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_entries_barrier_7_io_y_u; // @[package.scala 236:25]
  wire  tlb_entries_barrier_7_io_y_ae; // @[package.scala 236:25]
  wire  tlb_entries_barrier_7_io_y_sw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_7_io_y_sx; // @[package.scala 236:25]
  wire  tlb_entries_barrier_7_io_y_sr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_7_io_y_pw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_7_io_y_px; // @[package.scala 236:25]
  wire  tlb_entries_barrier_7_io_y_pr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_7_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_entries_barrier_7_io_y_pal; // @[package.scala 236:25]
  wire  tlb_entries_barrier_7_io_y_paa; // @[package.scala 236:25]
  wire  tlb_entries_barrier_7_io_y_eff; // @[package.scala 236:25]
  wire  tlb_entries_barrier_7_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_entries_barrier_8_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_entries_barrier_8_io_x_u; // @[package.scala 236:25]
  wire  tlb_entries_barrier_8_io_x_ae; // @[package.scala 236:25]
  wire  tlb_entries_barrier_8_io_x_sw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_8_io_x_sx; // @[package.scala 236:25]
  wire  tlb_entries_barrier_8_io_x_sr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_8_io_x_pw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_8_io_x_px; // @[package.scala 236:25]
  wire  tlb_entries_barrier_8_io_x_pr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_8_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_entries_barrier_8_io_x_pal; // @[package.scala 236:25]
  wire  tlb_entries_barrier_8_io_x_paa; // @[package.scala 236:25]
  wire  tlb_entries_barrier_8_io_x_eff; // @[package.scala 236:25]
  wire  tlb_entries_barrier_8_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_entries_barrier_8_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_entries_barrier_8_io_y_u; // @[package.scala 236:25]
  wire  tlb_entries_barrier_8_io_y_ae; // @[package.scala 236:25]
  wire  tlb_entries_barrier_8_io_y_sw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_8_io_y_sx; // @[package.scala 236:25]
  wire  tlb_entries_barrier_8_io_y_sr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_8_io_y_pw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_8_io_y_px; // @[package.scala 236:25]
  wire  tlb_entries_barrier_8_io_y_pr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_8_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_entries_barrier_8_io_y_pal; // @[package.scala 236:25]
  wire  tlb_entries_barrier_8_io_y_paa; // @[package.scala 236:25]
  wire  tlb_entries_barrier_8_io_y_eff; // @[package.scala 236:25]
  wire  tlb_entries_barrier_8_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_entries_barrier_9_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_entries_barrier_9_io_x_u; // @[package.scala 236:25]
  wire  tlb_entries_barrier_9_io_x_ae; // @[package.scala 236:25]
  wire  tlb_entries_barrier_9_io_x_sw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_9_io_x_sx; // @[package.scala 236:25]
  wire  tlb_entries_barrier_9_io_x_sr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_9_io_x_pw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_9_io_x_px; // @[package.scala 236:25]
  wire  tlb_entries_barrier_9_io_x_pr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_9_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_entries_barrier_9_io_x_pal; // @[package.scala 236:25]
  wire  tlb_entries_barrier_9_io_x_paa; // @[package.scala 236:25]
  wire  tlb_entries_barrier_9_io_x_eff; // @[package.scala 236:25]
  wire  tlb_entries_barrier_9_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_entries_barrier_9_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_entries_barrier_9_io_y_u; // @[package.scala 236:25]
  wire  tlb_entries_barrier_9_io_y_ae; // @[package.scala 236:25]
  wire  tlb_entries_barrier_9_io_y_sw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_9_io_y_sx; // @[package.scala 236:25]
  wire  tlb_entries_barrier_9_io_y_sr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_9_io_y_pw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_9_io_y_px; // @[package.scala 236:25]
  wire  tlb_entries_barrier_9_io_y_pr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_9_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_entries_barrier_9_io_y_pal; // @[package.scala 236:25]
  wire  tlb_entries_barrier_9_io_y_paa; // @[package.scala 236:25]
  wire  tlb_entries_barrier_9_io_y_eff; // @[package.scala 236:25]
  wire  tlb_entries_barrier_9_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_entries_barrier_10_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_entries_barrier_10_io_x_u; // @[package.scala 236:25]
  wire  tlb_entries_barrier_10_io_x_ae; // @[package.scala 236:25]
  wire  tlb_entries_barrier_10_io_x_sw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_10_io_x_sx; // @[package.scala 236:25]
  wire  tlb_entries_barrier_10_io_x_sr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_10_io_x_pw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_10_io_x_px; // @[package.scala 236:25]
  wire  tlb_entries_barrier_10_io_x_pr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_10_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_entries_barrier_10_io_x_pal; // @[package.scala 236:25]
  wire  tlb_entries_barrier_10_io_x_paa; // @[package.scala 236:25]
  wire  tlb_entries_barrier_10_io_x_eff; // @[package.scala 236:25]
  wire  tlb_entries_barrier_10_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_entries_barrier_10_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_entries_barrier_10_io_y_u; // @[package.scala 236:25]
  wire  tlb_entries_barrier_10_io_y_ae; // @[package.scala 236:25]
  wire  tlb_entries_barrier_10_io_y_sw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_10_io_y_sx; // @[package.scala 236:25]
  wire  tlb_entries_barrier_10_io_y_sr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_10_io_y_pw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_10_io_y_px; // @[package.scala 236:25]
  wire  tlb_entries_barrier_10_io_y_pr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_10_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_entries_barrier_10_io_y_pal; // @[package.scala 236:25]
  wire  tlb_entries_barrier_10_io_y_paa; // @[package.scala 236:25]
  wire  tlb_entries_barrier_10_io_y_eff; // @[package.scala 236:25]
  wire  tlb_entries_barrier_10_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_entries_barrier_11_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_entries_barrier_11_io_x_u; // @[package.scala 236:25]
  wire  tlb_entries_barrier_11_io_x_ae; // @[package.scala 236:25]
  wire  tlb_entries_barrier_11_io_x_sw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_11_io_x_sx; // @[package.scala 236:25]
  wire  tlb_entries_barrier_11_io_x_sr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_11_io_x_pw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_11_io_x_px; // @[package.scala 236:25]
  wire  tlb_entries_barrier_11_io_x_pr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_11_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_entries_barrier_11_io_x_pal; // @[package.scala 236:25]
  wire  tlb_entries_barrier_11_io_x_paa; // @[package.scala 236:25]
  wire  tlb_entries_barrier_11_io_x_eff; // @[package.scala 236:25]
  wire  tlb_entries_barrier_11_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_entries_barrier_11_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_entries_barrier_11_io_y_u; // @[package.scala 236:25]
  wire  tlb_entries_barrier_11_io_y_ae; // @[package.scala 236:25]
  wire  tlb_entries_barrier_11_io_y_sw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_11_io_y_sx; // @[package.scala 236:25]
  wire  tlb_entries_barrier_11_io_y_sr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_11_io_y_pw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_11_io_y_px; // @[package.scala 236:25]
  wire  tlb_entries_barrier_11_io_y_pr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_11_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_entries_barrier_11_io_y_pal; // @[package.scala 236:25]
  wire  tlb_entries_barrier_11_io_y_paa; // @[package.scala 236:25]
  wire  tlb_entries_barrier_11_io_y_eff; // @[package.scala 236:25]
  wire  tlb_entries_barrier_11_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_entries_barrier_12_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_entries_barrier_12_io_x_u; // @[package.scala 236:25]
  wire  tlb_entries_barrier_12_io_x_ae; // @[package.scala 236:25]
  wire  tlb_entries_barrier_12_io_x_sw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_12_io_x_sx; // @[package.scala 236:25]
  wire  tlb_entries_barrier_12_io_x_sr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_12_io_x_pw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_12_io_x_px; // @[package.scala 236:25]
  wire  tlb_entries_barrier_12_io_x_pr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_12_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_entries_barrier_12_io_x_pal; // @[package.scala 236:25]
  wire  tlb_entries_barrier_12_io_x_paa; // @[package.scala 236:25]
  wire  tlb_entries_barrier_12_io_x_eff; // @[package.scala 236:25]
  wire  tlb_entries_barrier_12_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_entries_barrier_12_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_entries_barrier_12_io_y_u; // @[package.scala 236:25]
  wire  tlb_entries_barrier_12_io_y_ae; // @[package.scala 236:25]
  wire  tlb_entries_barrier_12_io_y_sw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_12_io_y_sx; // @[package.scala 236:25]
  wire  tlb_entries_barrier_12_io_y_sr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_12_io_y_pw; // @[package.scala 236:25]
  wire  tlb_entries_barrier_12_io_y_px; // @[package.scala 236:25]
  wire  tlb_entries_barrier_12_io_y_pr; // @[package.scala 236:25]
  wire  tlb_entries_barrier_12_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_entries_barrier_12_io_y_pal; // @[package.scala 236:25]
  wire  tlb_entries_barrier_12_io_y_paa; // @[package.scala 236:25]
  wire  tlb_entries_barrier_12_io_y_eff; // @[package.scala 236:25]
  wire  tlb_entries_barrier_12_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_normal_entries_barrier_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_io_x_u; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_io_x_ae; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_io_x_sw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_io_x_sx; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_io_x_sr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_io_x_pw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_io_x_px; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_io_x_pr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_io_x_pal; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_io_x_paa; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_io_x_eff; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_normal_entries_barrier_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_io_y_u; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_io_y_ae; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_io_y_sw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_io_y_sx; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_io_y_sr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_io_y_pw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_io_y_px; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_io_y_pr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_io_y_pal; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_io_y_paa; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_io_y_eff; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_normal_entries_barrier_1_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_1_io_x_u; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_1_io_x_ae; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_1_io_x_sw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_1_io_x_sx; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_1_io_x_sr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_1_io_x_pw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_1_io_x_px; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_1_io_x_pr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_1_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_1_io_x_pal; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_1_io_x_paa; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_1_io_x_eff; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_1_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_normal_entries_barrier_1_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_1_io_y_u; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_1_io_y_ae; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_1_io_y_sw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_1_io_y_sx; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_1_io_y_sr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_1_io_y_pw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_1_io_y_px; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_1_io_y_pr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_1_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_1_io_y_pal; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_1_io_y_paa; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_1_io_y_eff; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_1_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_normal_entries_barrier_2_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_2_io_x_u; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_2_io_x_ae; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_2_io_x_sw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_2_io_x_sx; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_2_io_x_sr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_2_io_x_pw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_2_io_x_px; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_2_io_x_pr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_2_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_2_io_x_pal; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_2_io_x_paa; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_2_io_x_eff; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_2_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_normal_entries_barrier_2_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_2_io_y_u; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_2_io_y_ae; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_2_io_y_sw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_2_io_y_sx; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_2_io_y_sr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_2_io_y_pw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_2_io_y_px; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_2_io_y_pr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_2_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_2_io_y_pal; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_2_io_y_paa; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_2_io_y_eff; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_2_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_normal_entries_barrier_3_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_3_io_x_u; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_3_io_x_ae; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_3_io_x_sw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_3_io_x_sx; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_3_io_x_sr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_3_io_x_pw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_3_io_x_px; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_3_io_x_pr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_3_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_3_io_x_pal; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_3_io_x_paa; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_3_io_x_eff; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_3_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_normal_entries_barrier_3_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_3_io_y_u; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_3_io_y_ae; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_3_io_y_sw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_3_io_y_sx; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_3_io_y_sr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_3_io_y_pw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_3_io_y_px; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_3_io_y_pr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_3_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_3_io_y_pal; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_3_io_y_paa; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_3_io_y_eff; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_3_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_normal_entries_barrier_4_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_4_io_x_u; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_4_io_x_ae; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_4_io_x_sw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_4_io_x_sx; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_4_io_x_sr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_4_io_x_pw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_4_io_x_px; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_4_io_x_pr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_4_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_4_io_x_pal; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_4_io_x_paa; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_4_io_x_eff; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_4_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_normal_entries_barrier_4_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_4_io_y_u; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_4_io_y_ae; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_4_io_y_sw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_4_io_y_sx; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_4_io_y_sr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_4_io_y_pw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_4_io_y_px; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_4_io_y_pr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_4_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_4_io_y_pal; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_4_io_y_paa; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_4_io_y_eff; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_4_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_normal_entries_barrier_5_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_5_io_x_u; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_5_io_x_ae; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_5_io_x_sw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_5_io_x_sx; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_5_io_x_sr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_5_io_x_pw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_5_io_x_px; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_5_io_x_pr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_5_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_5_io_x_pal; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_5_io_x_paa; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_5_io_x_eff; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_5_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_normal_entries_barrier_5_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_5_io_y_u; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_5_io_y_ae; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_5_io_y_sw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_5_io_y_sx; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_5_io_y_sr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_5_io_y_pw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_5_io_y_px; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_5_io_y_pr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_5_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_5_io_y_pal; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_5_io_y_paa; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_5_io_y_eff; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_5_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_normal_entries_barrier_6_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_6_io_x_u; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_6_io_x_ae; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_6_io_x_sw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_6_io_x_sx; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_6_io_x_sr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_6_io_x_pw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_6_io_x_px; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_6_io_x_pr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_6_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_6_io_x_pal; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_6_io_x_paa; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_6_io_x_eff; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_6_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_normal_entries_barrier_6_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_6_io_y_u; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_6_io_y_ae; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_6_io_y_sw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_6_io_y_sx; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_6_io_y_sr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_6_io_y_pw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_6_io_y_px; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_6_io_y_pr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_6_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_6_io_y_pal; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_6_io_y_paa; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_6_io_y_eff; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_6_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_normal_entries_barrier_7_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_7_io_x_u; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_7_io_x_ae; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_7_io_x_sw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_7_io_x_sx; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_7_io_x_sr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_7_io_x_pw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_7_io_x_px; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_7_io_x_pr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_7_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_7_io_x_pal; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_7_io_x_paa; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_7_io_x_eff; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_7_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_normal_entries_barrier_7_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_7_io_y_u; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_7_io_y_ae; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_7_io_y_sw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_7_io_y_sx; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_7_io_y_sr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_7_io_y_pw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_7_io_y_px; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_7_io_y_pr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_7_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_7_io_y_pal; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_7_io_y_paa; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_7_io_y_eff; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_7_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_normal_entries_barrier_8_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_8_io_x_u; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_8_io_x_ae; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_8_io_x_sw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_8_io_x_sx; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_8_io_x_sr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_8_io_x_pw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_8_io_x_px; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_8_io_x_pr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_8_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_8_io_x_pal; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_8_io_x_paa; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_8_io_x_eff; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_8_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_normal_entries_barrier_8_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_8_io_y_u; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_8_io_y_ae; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_8_io_y_sw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_8_io_y_sx; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_8_io_y_sr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_8_io_y_pw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_8_io_y_px; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_8_io_y_pr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_8_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_8_io_y_pal; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_8_io_y_paa; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_8_io_y_eff; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_8_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_normal_entries_barrier_9_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_9_io_x_u; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_9_io_x_ae; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_9_io_x_sw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_9_io_x_sx; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_9_io_x_sr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_9_io_x_pw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_9_io_x_px; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_9_io_x_pr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_9_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_9_io_x_pal; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_9_io_x_paa; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_9_io_x_eff; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_9_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_normal_entries_barrier_9_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_9_io_y_u; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_9_io_y_ae; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_9_io_y_sw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_9_io_y_sx; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_9_io_y_sr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_9_io_y_pw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_9_io_y_px; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_9_io_y_pr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_9_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_9_io_y_pal; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_9_io_y_paa; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_9_io_y_eff; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_9_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_normal_entries_barrier_10_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_10_io_x_u; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_10_io_x_ae; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_10_io_x_sw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_10_io_x_sx; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_10_io_x_sr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_10_io_x_pw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_10_io_x_px; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_10_io_x_pr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_10_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_10_io_x_pal; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_10_io_x_paa; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_10_io_x_eff; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_10_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_normal_entries_barrier_10_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_10_io_y_u; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_10_io_y_ae; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_10_io_y_sw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_10_io_y_sx; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_10_io_y_sr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_10_io_y_pw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_10_io_y_px; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_10_io_y_pr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_10_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_10_io_y_pal; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_10_io_y_paa; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_10_io_y_eff; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_10_io_y_c; // @[package.scala 236:25]
  wire [19:0] tlb_normal_entries_barrier_11_io_x_ppn; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_11_io_x_u; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_11_io_x_ae; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_11_io_x_sw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_11_io_x_sx; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_11_io_x_sr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_11_io_x_pw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_11_io_x_px; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_11_io_x_pr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_11_io_x_ppp; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_11_io_x_pal; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_11_io_x_paa; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_11_io_x_eff; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_11_io_x_c; // @[package.scala 236:25]
  wire [19:0] tlb_normal_entries_barrier_11_io_y_ppn; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_11_io_y_u; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_11_io_y_ae; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_11_io_y_sw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_11_io_y_sx; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_11_io_y_sr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_11_io_y_pw; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_11_io_y_px; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_11_io_y_pr; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_11_io_y_ppp; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_11_io_y_pal; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_11_io_y_paa; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_11_io_y_eff; // @[package.scala 236:25]
  wire  tlb_normal_entries_barrier_11_io_y_c; // @[package.scala 236:25]
  reg [26:0] tlb_sectored_entries_0_tag; // @[TLB.scala 162:29]
  reg [34:0] tlb_sectored_entries_0_data_0; // @[TLB.scala 162:29]
  reg [34:0] tlb_sectored_entries_0_data_1; // @[TLB.scala 162:29]
  reg [34:0] tlb_sectored_entries_0_data_2; // @[TLB.scala 162:29]
  reg [34:0] tlb_sectored_entries_0_data_3; // @[TLB.scala 162:29]
  reg  tlb_sectored_entries_0_valid_0; // @[TLB.scala 162:29]
  reg  tlb_sectored_entries_0_valid_1; // @[TLB.scala 162:29]
  reg  tlb_sectored_entries_0_valid_2; // @[TLB.scala 162:29]
  reg  tlb_sectored_entries_0_valid_3; // @[TLB.scala 162:29]
  reg [26:0] tlb_sectored_entries_1_tag; // @[TLB.scala 162:29]
  reg [34:0] tlb_sectored_entries_1_data_0; // @[TLB.scala 162:29]
  reg [34:0] tlb_sectored_entries_1_data_1; // @[TLB.scala 162:29]
  reg [34:0] tlb_sectored_entries_1_data_2; // @[TLB.scala 162:29]
  reg [34:0] tlb_sectored_entries_1_data_3; // @[TLB.scala 162:29]
  reg  tlb_sectored_entries_1_valid_0; // @[TLB.scala 162:29]
  reg  tlb_sectored_entries_1_valid_1; // @[TLB.scala 162:29]
  reg  tlb_sectored_entries_1_valid_2; // @[TLB.scala 162:29]
  reg  tlb_sectored_entries_1_valid_3; // @[TLB.scala 162:29]
  reg [26:0] tlb_sectored_entries_2_tag; // @[TLB.scala 162:29]
  reg [34:0] tlb_sectored_entries_2_data_0; // @[TLB.scala 162:29]
  reg [34:0] tlb_sectored_entries_2_data_1; // @[TLB.scala 162:29]
  reg [34:0] tlb_sectored_entries_2_data_2; // @[TLB.scala 162:29]
  reg [34:0] tlb_sectored_entries_2_data_3; // @[TLB.scala 162:29]
  reg  tlb_sectored_entries_2_valid_0; // @[TLB.scala 162:29]
  reg  tlb_sectored_entries_2_valid_1; // @[TLB.scala 162:29]
  reg  tlb_sectored_entries_2_valid_2; // @[TLB.scala 162:29]
  reg  tlb_sectored_entries_2_valid_3; // @[TLB.scala 162:29]
  reg [26:0] tlb_sectored_entries_3_tag; // @[TLB.scala 162:29]
  reg [34:0] tlb_sectored_entries_3_data_0; // @[TLB.scala 162:29]
  reg [34:0] tlb_sectored_entries_3_data_1; // @[TLB.scala 162:29]
  reg [34:0] tlb_sectored_entries_3_data_2; // @[TLB.scala 162:29]
  reg [34:0] tlb_sectored_entries_3_data_3; // @[TLB.scala 162:29]
  reg  tlb_sectored_entries_3_valid_0; // @[TLB.scala 162:29]
  reg  tlb_sectored_entries_3_valid_1; // @[TLB.scala 162:29]
  reg  tlb_sectored_entries_3_valid_2; // @[TLB.scala 162:29]
  reg  tlb_sectored_entries_3_valid_3; // @[TLB.scala 162:29]
  reg [26:0] tlb_sectored_entries_4_tag; // @[TLB.scala 162:29]
  reg [34:0] tlb_sectored_entries_4_data_0; // @[TLB.scala 162:29]
  reg [34:0] tlb_sectored_entries_4_data_1; // @[TLB.scala 162:29]
  reg [34:0] tlb_sectored_entries_4_data_2; // @[TLB.scala 162:29]
  reg [34:0] tlb_sectored_entries_4_data_3; // @[TLB.scala 162:29]
  reg  tlb_sectored_entries_4_valid_0; // @[TLB.scala 162:29]
  reg  tlb_sectored_entries_4_valid_1; // @[TLB.scala 162:29]
  reg  tlb_sectored_entries_4_valid_2; // @[TLB.scala 162:29]
  reg  tlb_sectored_entries_4_valid_3; // @[TLB.scala 162:29]
  reg [26:0] tlb_sectored_entries_5_tag; // @[TLB.scala 162:29]
  reg [34:0] tlb_sectored_entries_5_data_0; // @[TLB.scala 162:29]
  reg [34:0] tlb_sectored_entries_5_data_1; // @[TLB.scala 162:29]
  reg [34:0] tlb_sectored_entries_5_data_2; // @[TLB.scala 162:29]
  reg [34:0] tlb_sectored_entries_5_data_3; // @[TLB.scala 162:29]
  reg  tlb_sectored_entries_5_valid_0; // @[TLB.scala 162:29]
  reg  tlb_sectored_entries_5_valid_1; // @[TLB.scala 162:29]
  reg  tlb_sectored_entries_5_valid_2; // @[TLB.scala 162:29]
  reg  tlb_sectored_entries_5_valid_3; // @[TLB.scala 162:29]
  reg [26:0] tlb_sectored_entries_6_tag; // @[TLB.scala 162:29]
  reg [34:0] tlb_sectored_entries_6_data_0; // @[TLB.scala 162:29]
  reg [34:0] tlb_sectored_entries_6_data_1; // @[TLB.scala 162:29]
  reg [34:0] tlb_sectored_entries_6_data_2; // @[TLB.scala 162:29]
  reg [34:0] tlb_sectored_entries_6_data_3; // @[TLB.scala 162:29]
  reg  tlb_sectored_entries_6_valid_0; // @[TLB.scala 162:29]
  reg  tlb_sectored_entries_6_valid_1; // @[TLB.scala 162:29]
  reg  tlb_sectored_entries_6_valid_2; // @[TLB.scala 162:29]
  reg  tlb_sectored_entries_6_valid_3; // @[TLB.scala 162:29]
  reg [26:0] tlb_sectored_entries_7_tag; // @[TLB.scala 162:29]
  reg [34:0] tlb_sectored_entries_7_data_0; // @[TLB.scala 162:29]
  reg [34:0] tlb_sectored_entries_7_data_1; // @[TLB.scala 162:29]
  reg [34:0] tlb_sectored_entries_7_data_2; // @[TLB.scala 162:29]
  reg [34:0] tlb_sectored_entries_7_data_3; // @[TLB.scala 162:29]
  reg  tlb_sectored_entries_7_valid_0; // @[TLB.scala 162:29]
  reg  tlb_sectored_entries_7_valid_1; // @[TLB.scala 162:29]
  reg  tlb_sectored_entries_7_valid_2; // @[TLB.scala 162:29]
  reg  tlb_sectored_entries_7_valid_3; // @[TLB.scala 162:29]
  reg [1:0] tlb_superpage_entries_0_level; // @[TLB.scala 163:30]
  reg [26:0] tlb_superpage_entries_0_tag; // @[TLB.scala 163:30]
  reg [34:0] tlb_superpage_entries_0_data_0; // @[TLB.scala 163:30]
  reg  tlb_superpage_entries_0_valid_0; // @[TLB.scala 163:30]
  reg [1:0] tlb_superpage_entries_1_level; // @[TLB.scala 163:30]
  reg [26:0] tlb_superpage_entries_1_tag; // @[TLB.scala 163:30]
  reg [34:0] tlb_superpage_entries_1_data_0; // @[TLB.scala 163:30]
  reg  tlb_superpage_entries_1_valid_0; // @[TLB.scala 163:30]
  reg [1:0] tlb_superpage_entries_2_level; // @[TLB.scala 163:30]
  reg [26:0] tlb_superpage_entries_2_tag; // @[TLB.scala 163:30]
  reg [34:0] tlb_superpage_entries_2_data_0; // @[TLB.scala 163:30]
  reg  tlb_superpage_entries_2_valid_0; // @[TLB.scala 163:30]
  reg [1:0] tlb_superpage_entries_3_level; // @[TLB.scala 163:30]
  reg [26:0] tlb_superpage_entries_3_tag; // @[TLB.scala 163:30]
  reg [34:0] tlb_superpage_entries_3_data_0; // @[TLB.scala 163:30]
  reg  tlb_superpage_entries_3_valid_0; // @[TLB.scala 163:30]
  reg [1:0] tlb_special_entry_level; // @[TLB.scala 164:56]
  reg [26:0] tlb_special_entry_tag; // @[TLB.scala 164:56]
  reg [34:0] tlb_special_entry_data_0; // @[TLB.scala 164:56]
  reg  tlb_special_entry_valid_0; // @[TLB.scala 164:56]
  reg [1:0] tlb_state; // @[TLB.scala 169:18]
  reg [26:0] tlb_r_refill_tag; // @[TLB.scala 170:25]
  reg [1:0] tlb_r_superpage_repl_addr; // @[TLB.scala 171:34]
  reg [2:0] tlb_r_sectored_repl_addr; // @[TLB.scala 172:33]
  reg [2:0] tlb_r_sectored_hit_addr; // @[TLB.scala 173:32]
  reg  tlb_r_sectored_hit; // @[TLB.scala 174:27]
  wire  tlb_priv_s = tlb_io_ptw_status_dprv[0]; // @[TLB.scala 177:20]
  wire  tlb_priv_uses_vm = tlb_io_ptw_status_dprv <= 2'h1; // @[TLB.scala 178:27]
  wire  tlb__vm_enabled_T = tlb_io_ptw_ptbr_mode[3]; // @[TLB.scala 179:53]
  wire  tlb__vm_enabled_T_2 = tlb__vm_enabled_T & tlb_priv_uses_vm; // @[TLB.scala 179:83]
  wire  tlb__vm_enabled_T_3 = ~tlb_io_req_bits_passthrough; // @[TLB.scala 179:102]
  wire  tlb_vm_enabled = tlb__vm_enabled_T_2 & tlb__vm_enabled_T_3; // @[TLB.scala 179:99]
  wire [26:0] tlb_vpn = tlb_io_req_bits_vaddr[38:12]; // @[TLB.scala 182:30]
  wire [19:0] tlb_refill_ppn = tlb_io_ptw_resp_bits_pte_ppn[19:0]; // @[TLB.scala 183:44]
  wire  tlb__invalidate_refill_T = tlb_state == 2'h1; // @[package.scala 15:47]
  wire  tlb__invalidate_refill_T_1 = tlb_state == 2'h3; // @[package.scala 15:47]
  wire  tlb__invalidate_refill_T_2 = tlb__invalidate_refill_T | tlb__invalidate_refill_T_1; // @[package.scala 64:59]
  wire  tlb_invalidate_refill = tlb__invalidate_refill_T_2 | tlb_io_sfence_valid; // @[TLB.scala 185:88]
  wire  tlb__mpu_ppn_data_T_13 = tlb_special_entry_data_0[13]; // @[TLB.scala 86:77]
  wire [1:0] tlb_mpu_ppn_right = tlb_mpu_ppn_data_barrier_io_y_ppn[19:18]; // @[TLB.scala 106:26]
  wire  tlb__mpu_ppn_ignore_T = tlb_special_entry_level < 2'h1; // @[TLB.scala 108:28]
  wire [26:0] tlb__mpu_ppn_T_1 = tlb__mpu_ppn_ignore_T ? tlb_vpn : 27'h0; // @[TLB.scala 109:28]
  wire [26:0] _GEN_347 = {{7'd0}, tlb_mpu_ppn_data_barrier_io_y_ppn}; // @[TLB.scala 109:47]
  wire [26:0] tlb__mpu_ppn_T_2 = tlb__mpu_ppn_T_1 | _GEN_347; // @[TLB.scala 109:47]
  wire [8:0] tlb_mpu_ppn_left = tlb__mpu_ppn_T_2[17:9]; // @[TLB.scala 109:58]
  wire  tlb__mpu_ppn_ignore_T_1 = tlb_special_entry_level < 2'h2; // @[TLB.scala 108:28]
  wire [26:0] tlb__mpu_ppn_T_3 = tlb__mpu_ppn_ignore_T_1 ? tlb_vpn : 27'h0; // @[TLB.scala 109:28]
  wire [26:0] tlb__mpu_ppn_T_4 = tlb__mpu_ppn_T_3 | _GEN_347; // @[TLB.scala 109:47]
  wire [8:0] tlb_mpu_ppn_left_1 = tlb__mpu_ppn_T_4[8:0]; // @[TLB.scala 109:58]
  wire [19:0] tlb__mpu_ppn_T_5 = {tlb_mpu_ppn_right,tlb_mpu_ppn_left,tlb_mpu_ppn_left_1}; // @[Cat.scala 29:58]
  wire [27:0] tlb__mpu_ppn_T_6 = tlb_io_req_bits_vaddr[39:12]; // @[TLB.scala 187:123]
  wire [27:0] tlb__mpu_ppn_T_7 = tlb_vm_enabled ? {{8'd0}, tlb__mpu_ppn_T_5} : tlb__mpu_ppn_T_6; // @[TLB.scala 187:20]
  wire [27:0] tlb_mpu_ppn = tlb_io_ptw_resp_valid ? {{8'd0}, tlb_refill_ppn} : tlb__mpu_ppn_T_7; // @[TLB.scala 186:20]
  wire [11:0] tlb_mpu_physaddr_left = tlb_io_req_bits_vaddr[11:0]; // @[TLB.scala 188:52]
  wire [39:0] tlb_mpu_physaddr = {tlb_mpu_ppn,tlb_mpu_physaddr_left}; // @[Cat.scala 29:58]
  wire  tlb__mpu_priv_T = tlb_io_ptw_resp_valid | tlb_io_req_bits_passthrough; // @[TLB.scala 189:56]
  wire [2:0] tlb__mpu_priv_T_2 = {tlb_io_ptw_status_debug,tlb_io_ptw_status_dprv}; // @[Cat.scala 29:58]
  wire [2:0] tlb_mpu_priv = tlb__mpu_priv_T ? 3'h1 : tlb__mpu_priv_T_2; // @[TLB.scala 189:27]
  wire [39:0] tlb__legal_address_T = tlb_mpu_physaddr ^ 40'h3000; // @[Parameters.scala 138:31]
  wire [40:0] tlb__legal_address_T_1 = {1'b0,$signed(tlb__legal_address_T)}; // @[Parameters.scala 138:49]
  wire [40:0] tlb__legal_address_T_3 = $signed(tlb__legal_address_T_1) & -41'sh1000; // @[Parameters.scala 138:52]
  wire  tlb__legal_address_T_4 = $signed(tlb__legal_address_T_3) == 41'sh0; // @[Parameters.scala 138:67]
  wire [39:0] tlb__legal_address_T_5 = tlb_mpu_physaddr ^ 40'hc000000; // @[Parameters.scala 138:31]
  wire [40:0] tlb__legal_address_T_6 = {1'b0,$signed(tlb__legal_address_T_5)}; // @[Parameters.scala 138:49]
  wire [40:0] tlb__legal_address_T_8 = $signed(tlb__legal_address_T_6) & -41'sh4000000; // @[Parameters.scala 138:52]
  wire  tlb__legal_address_T_9 = $signed(tlb__legal_address_T_8) == 41'sh0; // @[Parameters.scala 138:67]
  wire [39:0] tlb__legal_address_T_10 = tlb_mpu_physaddr ^ 40'h2000000; // @[Parameters.scala 138:31]
  wire [40:0] tlb__legal_address_T_11 = {1'b0,$signed(tlb__legal_address_T_10)}; // @[Parameters.scala 138:49]
  wire [40:0] tlb__legal_address_T_13 = $signed(tlb__legal_address_T_11) & -41'sh10000; // @[Parameters.scala 138:52]
  wire  tlb__legal_address_T_14 = $signed(tlb__legal_address_T_13) == 41'sh0; // @[Parameters.scala 138:67]
  wire [40:0] tlb__legal_address_T_16 = {1'b0,$signed(tlb_mpu_physaddr)}; // @[Parameters.scala 138:49]
  wire [40:0] tlb__legal_address_T_18 = $signed(tlb__legal_address_T_16) & -41'sh1000; // @[Parameters.scala 138:52]
  wire  tlb__legal_address_T_19 = $signed(tlb__legal_address_T_18) == 41'sh0; // @[Parameters.scala 138:67]
  wire [39:0] tlb__legal_address_T_20 = tlb_mpu_physaddr ^ 40'h10000; // @[Parameters.scala 138:31]
  wire [40:0] tlb__legal_address_T_21 = {1'b0,$signed(tlb__legal_address_T_20)}; // @[Parameters.scala 138:49]
  wire [40:0] tlb__legal_address_T_23 = $signed(tlb__legal_address_T_21) & -41'sh10000; // @[Parameters.scala 138:52]
  wire  tlb__legal_address_T_24 = $signed(tlb__legal_address_T_23) == 41'sh0; // @[Parameters.scala 138:67]
  wire [39:0] tlb__legal_address_T_25 = tlb_mpu_physaddr ^ 40'h80000000; // @[Parameters.scala 138:31]
  wire [40:0] tlb__legal_address_T_26 = {1'b0,$signed(tlb__legal_address_T_25)}; // @[Parameters.scala 138:49]
  wire [40:0] tlb__legal_address_T_28 = $signed(tlb__legal_address_T_26) & -41'sh10000000; // @[Parameters.scala 138:52]
  wire  tlb__legal_address_T_29 = $signed(tlb__legal_address_T_28) == 41'sh0; // @[Parameters.scala 138:67]
  wire [39:0] tlb__legal_address_T_30 = tlb_mpu_physaddr ^ 40'h60000000; // @[Parameters.scala 138:31]
  wire [40:0] tlb__legal_address_T_31 = {1'b0,$signed(tlb__legal_address_T_30)}; // @[Parameters.scala 138:49]
  wire [40:0] tlb__legal_address_T_33 = $signed(tlb__legal_address_T_31) & -41'sh20000000; // @[Parameters.scala 138:52]
  wire  tlb__legal_address_T_34 = $signed(tlb__legal_address_T_33) == 41'sh0; // @[Parameters.scala 138:67]
  wire  tlb__legal_address_T_35 = tlb__legal_address_T_4 | tlb__legal_address_T_9; // @[TLB.scala 195:67]
  wire  tlb__legal_address_T_36 = tlb__legal_address_T_35 | tlb__legal_address_T_14; // @[TLB.scala 195:67]
  wire  tlb__legal_address_T_37 = tlb__legal_address_T_36 | tlb__legal_address_T_19; // @[TLB.scala 195:67]
  wire  tlb__legal_address_T_38 = tlb__legal_address_T_37 | tlb__legal_address_T_24; // @[TLB.scala 195:67]
  wire  tlb__legal_address_T_39 = tlb__legal_address_T_38 | tlb__legal_address_T_29; // @[TLB.scala 195:67]
  wire  tlb_legal_address = tlb__legal_address_T_39 | tlb__legal_address_T_34; // @[TLB.scala 195:67]
  wire [40:0] tlb__cacheable_T_8 = $signed(tlb__legal_address_T_26) & 41'sh80000000; // @[Parameters.scala 138:52]
  wire  tlb__cacheable_T_9 = $signed(tlb__cacheable_T_8) == 41'sh0; // @[Parameters.scala 138:67]
  wire  tlb__cacheable_T_13 = tlb_legal_address & tlb__cacheable_T_9; // @[TLB.scala 197:19]
  wire [39:0] tlb__homogeneous_T_54 = tlb_mpu_physaddr ^ 40'h8000000; // @[Parameters.scala 138:31]
  wire [40:0] tlb__homogeneous_T_55 = {1'b0,$signed(tlb__homogeneous_T_54)}; // @[Parameters.scala 138:49]
  wire [40:0] tlb__homogeneous_T_57 = $signed(tlb__homogeneous_T_55) & 41'shc8000000; // @[Parameters.scala 138:52]
  wire  tlb__homogeneous_T_58 = $signed(tlb__homogeneous_T_57) == 41'sh0; // @[Parameters.scala 138:67]
  wire [40:0] tlb__homogeneous_T_71 = $signed(tlb__legal_address_T_16) & 41'shc8010000; // @[Parameters.scala 138:52]
  wire  tlb__homogeneous_T_72 = $signed(tlb__homogeneous_T_71) == 41'sh0; // @[Parameters.scala 138:67]
  wire  tlb__homogeneous_T_79 = tlb__homogeneous_T_72 | tlb__homogeneous_T_58; // @[TLBPermissions.scala 82:66]
  wire  tlb__deny_access_to_debug_T = tlb_mpu_priv <= 3'h3; // @[TLB.scala 200:39]
  wire  tlb_deny_access_to_debug = tlb__deny_access_to_debug_T & tlb__legal_address_T_19; // @[TLB.scala 200:48]
  wire  tlb__prot_r_T_6 = ~tlb_deny_access_to_debug; // @[TLB.scala 201:44]
  wire  tlb__prot_r_T_7 = tlb_legal_address & tlb__prot_r_T_6; // @[TLB.scala 201:41]
  wire  tlb_prot_r = tlb__prot_r_T_7 & tlb_pmp_io_r; // @[TLB.scala 201:66]
  wire [39:0] tlb__prot_w_T_10 = tlb_mpu_physaddr ^ 40'h40000000; // @[Parameters.scala 138:31]
  wire [40:0] tlb__prot_w_T_11 = {1'b0,$signed(tlb__prot_w_T_10)}; // @[Parameters.scala 138:49]
  wire [40:0] tlb__prot_w_T_13 = $signed(tlb__prot_w_T_11) & 41'shc0000000; // @[Parameters.scala 138:52]
  wire  tlb__prot_w_T_14 = $signed(tlb__prot_w_T_13) == 41'sh0; // @[Parameters.scala 138:67]
  wire [40:0] tlb__prot_w_T_18 = $signed(tlb__legal_address_T_26) & 41'shc0000000; // @[Parameters.scala 138:52]
  wire  tlb__prot_w_T_19 = $signed(tlb__prot_w_T_18) == 41'sh0; // @[Parameters.scala 138:67]
  wire  tlb__prot_w_T_21 = tlb__homogeneous_T_79 | tlb__prot_w_T_14; // @[Parameters.scala 616:89]
  wire  tlb__prot_w_T_22 = tlb__prot_w_T_21 | tlb__prot_w_T_19; // @[Parameters.scala 616:89]
  wire  tlb__prot_w_T_31 = tlb_legal_address & tlb__prot_w_T_22; // @[TLB.scala 197:19]
  wire  tlb__prot_w_T_33 = tlb__prot_w_T_31 & tlb__prot_r_T_6; // @[TLB.scala 202:45]
  wire  tlb_prot_w = tlb__prot_w_T_33 & tlb_pmp_io_w; // @[TLB.scala 202:70]
  wire  tlb_prot_al = tlb_legal_address & tlb__homogeneous_T_79; // @[TLB.scala 197:19]
  wire [40:0] tlb__prot_x_T_3 = $signed(tlb__legal_address_T_16) & 41'shca000000; // @[Parameters.scala 138:52]
  wire  tlb__prot_x_T_4 = $signed(tlb__prot_x_T_3) == 41'sh0; // @[Parameters.scala 138:67]
  wire  tlb__prot_x_T_15 = tlb__prot_x_T_4 | tlb__prot_w_T_14; // @[Parameters.scala 616:89]
  wire  tlb__prot_x_T_16 = tlb__prot_x_T_15 | tlb__prot_w_T_19; // @[Parameters.scala 616:89]
  wire  tlb__prot_x_T_31 = tlb_legal_address & tlb__prot_x_T_16; // @[TLB.scala 197:19]
  wire  tlb__prot_x_T_33 = tlb__prot_x_T_31 & tlb__prot_r_T_6; // @[TLB.scala 206:40]
  wire  tlb_prot_x = tlb__prot_x_T_33 & tlb_pmp_io_x; // @[TLB.scala 206:65]
  wire [40:0] tlb__prot_eff_T_20 = $signed(tlb__legal_address_T_16) & 41'shca012000; // @[Parameters.scala 138:52]
  wire  tlb__prot_eff_T_21 = $signed(tlb__prot_eff_T_20) == 41'sh0; // @[Parameters.scala 138:67]
  wire [40:0] tlb__prot_eff_T_25 = $signed(tlb__legal_address_T_11) & 41'shca010000; // @[Parameters.scala 138:52]
  wire  tlb__prot_eff_T_26 = $signed(tlb__prot_eff_T_25) == 41'sh0; // @[Parameters.scala 138:67]
  wire  tlb__prot_eff_T_37 = tlb__prot_eff_T_21 | tlb__prot_eff_T_26; // @[Parameters.scala 616:89]
  wire  tlb__prot_eff_T_38 = tlb__prot_eff_T_37 | tlb__homogeneous_T_58; // @[Parameters.scala 616:89]
  wire  tlb__prot_eff_T_39 = tlb__prot_eff_T_38 | tlb__prot_w_T_14; // @[Parameters.scala 616:89]
  wire  tlb_prot_eff = tlb_legal_address & tlb__prot_eff_T_39; // @[TLB.scala 197:19]
  wire  tlb__sector_hits_T = tlb_sectored_entries_0_valid_0 | tlb_sectored_entries_0_valid_1; // @[package.scala 64:59]
  wire  tlb__sector_hits_T_1 = tlb__sector_hits_T | tlb_sectored_entries_0_valid_2; // @[package.scala 64:59]
  wire  tlb__sector_hits_T_2 = tlb__sector_hits_T_1 | tlb_sectored_entries_0_valid_3; // @[package.scala 64:59]
  wire [26:0] tlb__sector_hits_T_3 = tlb_sectored_entries_0_tag ^ tlb_vpn; // @[TLB.scala 88:41]
  wire [24:0] tlb__sector_hits_T_4 = tlb__sector_hits_T_3[26:2]; // @[TLB.scala 88:48]
  wire  tlb__sector_hits_T_5 = tlb__sector_hits_T_4 == 25'h0; // @[TLB.scala 88:66]
  wire  tlb_sector_hits_0 = tlb__sector_hits_T_2 & tlb__sector_hits_T_5; // @[TLB.scala 87:40]
  wire  tlb__sector_hits_T_6 = tlb_sectored_entries_1_valid_0 | tlb_sectored_entries_1_valid_1; // @[package.scala 64:59]
  wire  tlb__sector_hits_T_7 = tlb__sector_hits_T_6 | tlb_sectored_entries_1_valid_2; // @[package.scala 64:59]
  wire  tlb__sector_hits_T_8 = tlb__sector_hits_T_7 | tlb_sectored_entries_1_valid_3; // @[package.scala 64:59]
  wire [26:0] tlb__sector_hits_T_9 = tlb_sectored_entries_1_tag ^ tlb_vpn; // @[TLB.scala 88:41]
  wire [24:0] tlb__sector_hits_T_10 = tlb__sector_hits_T_9[26:2]; // @[TLB.scala 88:48]
  wire  tlb__sector_hits_T_11 = tlb__sector_hits_T_10 == 25'h0; // @[TLB.scala 88:66]
  wire  tlb_sector_hits_1 = tlb__sector_hits_T_8 & tlb__sector_hits_T_11; // @[TLB.scala 87:40]
  wire  tlb__sector_hits_T_12 = tlb_sectored_entries_2_valid_0 | tlb_sectored_entries_2_valid_1; // @[package.scala 64:59]
  wire  tlb__sector_hits_T_13 = tlb__sector_hits_T_12 | tlb_sectored_entries_2_valid_2; // @[package.scala 64:59]
  wire  tlb__sector_hits_T_14 = tlb__sector_hits_T_13 | tlb_sectored_entries_2_valid_3; // @[package.scala 64:59]
  wire [26:0] tlb__sector_hits_T_15 = tlb_sectored_entries_2_tag ^ tlb_vpn; // @[TLB.scala 88:41]
  wire [24:0] tlb__sector_hits_T_16 = tlb__sector_hits_T_15[26:2]; // @[TLB.scala 88:48]
  wire  tlb__sector_hits_T_17 = tlb__sector_hits_T_16 == 25'h0; // @[TLB.scala 88:66]
  wire  tlb_sector_hits_2 = tlb__sector_hits_T_14 & tlb__sector_hits_T_17; // @[TLB.scala 87:40]
  wire  tlb__sector_hits_T_18 = tlb_sectored_entries_3_valid_0 | tlb_sectored_entries_3_valid_1; // @[package.scala 64:59]
  wire  tlb__sector_hits_T_19 = tlb__sector_hits_T_18 | tlb_sectored_entries_3_valid_2; // @[package.scala 64:59]
  wire  tlb__sector_hits_T_20 = tlb__sector_hits_T_19 | tlb_sectored_entries_3_valid_3; // @[package.scala 64:59]
  wire [26:0] tlb__sector_hits_T_21 = tlb_sectored_entries_3_tag ^ tlb_vpn; // @[TLB.scala 88:41]
  wire [24:0] tlb__sector_hits_T_22 = tlb__sector_hits_T_21[26:2]; // @[TLB.scala 88:48]
  wire  tlb__sector_hits_T_23 = tlb__sector_hits_T_22 == 25'h0; // @[TLB.scala 88:66]
  wire  tlb_sector_hits_3 = tlb__sector_hits_T_20 & tlb__sector_hits_T_23; // @[TLB.scala 87:40]
  wire  tlb__sector_hits_T_24 = tlb_sectored_entries_4_valid_0 | tlb_sectored_entries_4_valid_1; // @[package.scala 64:59]
  wire  tlb__sector_hits_T_25 = tlb__sector_hits_T_24 | tlb_sectored_entries_4_valid_2; // @[package.scala 64:59]
  wire  tlb__sector_hits_T_26 = tlb__sector_hits_T_25 | tlb_sectored_entries_4_valid_3; // @[package.scala 64:59]
  wire [26:0] tlb__sector_hits_T_27 = tlb_sectored_entries_4_tag ^ tlb_vpn; // @[TLB.scala 88:41]
  wire [24:0] tlb__sector_hits_T_28 = tlb__sector_hits_T_27[26:2]; // @[TLB.scala 88:48]
  wire  tlb__sector_hits_T_29 = tlb__sector_hits_T_28 == 25'h0; // @[TLB.scala 88:66]
  wire  tlb_sector_hits_4 = tlb__sector_hits_T_26 & tlb__sector_hits_T_29; // @[TLB.scala 87:40]
  wire  tlb__sector_hits_T_30 = tlb_sectored_entries_5_valid_0 | tlb_sectored_entries_5_valid_1; // @[package.scala 64:59]
  wire  tlb__sector_hits_T_31 = tlb__sector_hits_T_30 | tlb_sectored_entries_5_valid_2; // @[package.scala 64:59]
  wire  tlb__sector_hits_T_32 = tlb__sector_hits_T_31 | tlb_sectored_entries_5_valid_3; // @[package.scala 64:59]
  wire [26:0] tlb__sector_hits_T_33 = tlb_sectored_entries_5_tag ^ tlb_vpn; // @[TLB.scala 88:41]
  wire [24:0] tlb__sector_hits_T_34 = tlb__sector_hits_T_33[26:2]; // @[TLB.scala 88:48]
  wire  tlb__sector_hits_T_35 = tlb__sector_hits_T_34 == 25'h0; // @[TLB.scala 88:66]
  wire  tlb_sector_hits_5 = tlb__sector_hits_T_32 & tlb__sector_hits_T_35; // @[TLB.scala 87:40]
  wire  tlb__sector_hits_T_36 = tlb_sectored_entries_6_valid_0 | tlb_sectored_entries_6_valid_1; // @[package.scala 64:59]
  wire  tlb__sector_hits_T_37 = tlb__sector_hits_T_36 | tlb_sectored_entries_6_valid_2; // @[package.scala 64:59]
  wire  tlb__sector_hits_T_38 = tlb__sector_hits_T_37 | tlb_sectored_entries_6_valid_3; // @[package.scala 64:59]
  wire [26:0] tlb__sector_hits_T_39 = tlb_sectored_entries_6_tag ^ tlb_vpn; // @[TLB.scala 88:41]
  wire [24:0] tlb__sector_hits_T_40 = tlb__sector_hits_T_39[26:2]; // @[TLB.scala 88:48]
  wire  tlb__sector_hits_T_41 = tlb__sector_hits_T_40 == 25'h0; // @[TLB.scala 88:66]
  wire  tlb_sector_hits_6 = tlb__sector_hits_T_38 & tlb__sector_hits_T_41; // @[TLB.scala 87:40]
  wire  tlb__sector_hits_T_42 = tlb_sectored_entries_7_valid_0 | tlb_sectored_entries_7_valid_1; // @[package.scala 64:59]
  wire  tlb__sector_hits_T_43 = tlb__sector_hits_T_42 | tlb_sectored_entries_7_valid_2; // @[package.scala 64:59]
  wire  tlb__sector_hits_T_44 = tlb__sector_hits_T_43 | tlb_sectored_entries_7_valid_3; // @[package.scala 64:59]
  wire [26:0] tlb__sector_hits_T_45 = tlb_sectored_entries_7_tag ^ tlb_vpn; // @[TLB.scala 88:41]
  wire [24:0] tlb__sector_hits_T_46 = tlb__sector_hits_T_45[26:2]; // @[TLB.scala 88:48]
  wire  tlb__sector_hits_T_47 = tlb__sector_hits_T_46 == 25'h0; // @[TLB.scala 88:66]
  wire  tlb_sector_hits_7 = tlb__sector_hits_T_44 & tlb__sector_hits_T_47; // @[TLB.scala 87:40]
  wire [8:0] tlb__superpage_hits_T = tlb_superpage_entries_0_tag[26:18]; // @[TLB.scala 95:46]
  wire [8:0] tlb__superpage_hits_T_1 = tlb_vpn[26:18]; // @[TLB.scala 95:84]
  wire  tlb__superpage_hits_T_2 = tlb__superpage_hits_T == tlb__superpage_hits_T_1; // @[TLB.scala 95:77]
  wire  tlb__superpage_hits_T_4 = tlb_superpage_entries_0_valid_0 & tlb__superpage_hits_T_2; // @[TLB.scala 95:29]
  wire  tlb__superpage_hits_ignore_T_1 = tlb_superpage_entries_0_level < 2'h1; // @[TLB.scala 94:28]
  wire [8:0] tlb__superpage_hits_T_5 = tlb_superpage_entries_0_tag[17:9]; // @[TLB.scala 95:46]
  wire [8:0] tlb__superpage_hits_T_6 = tlb_vpn[17:9]; // @[TLB.scala 95:84]
  wire  tlb__superpage_hits_T_7 = tlb__superpage_hits_T_5 == tlb__superpage_hits_T_6; // @[TLB.scala 95:77]
  wire  tlb__superpage_hits_T_8 = tlb__superpage_hits_ignore_T_1 | tlb__superpage_hits_T_7; // @[TLB.scala 95:40]
  wire  tlb__superpage_hits_T_9 = tlb__superpage_hits_T_4 & tlb__superpage_hits_T_8; // @[TLB.scala 95:29]
  wire [8:0] tlb__superpage_hits_T_11 = tlb_vpn[8:0]; // @[TLB.scala 95:84]
  wire [8:0] tlb__superpage_hits_T_14 = tlb_superpage_entries_1_tag[26:18]; // @[TLB.scala 95:46]
  wire  tlb__superpage_hits_T_16 = tlb__superpage_hits_T_14 == tlb__superpage_hits_T_1; // @[TLB.scala 95:77]
  wire  tlb__superpage_hits_T_18 = tlb_superpage_entries_1_valid_0 & tlb__superpage_hits_T_16; // @[TLB.scala 95:29]
  wire  tlb__superpage_hits_ignore_T_4 = tlb_superpage_entries_1_level < 2'h1; // @[TLB.scala 94:28]
  wire [8:0] tlb__superpage_hits_T_19 = tlb_superpage_entries_1_tag[17:9]; // @[TLB.scala 95:46]
  wire  tlb__superpage_hits_T_21 = tlb__superpage_hits_T_19 == tlb__superpage_hits_T_6; // @[TLB.scala 95:77]
  wire  tlb__superpage_hits_T_22 = tlb__superpage_hits_ignore_T_4 | tlb__superpage_hits_T_21; // @[TLB.scala 95:40]
  wire  tlb__superpage_hits_T_23 = tlb__superpage_hits_T_18 & tlb__superpage_hits_T_22; // @[TLB.scala 95:29]
  wire [8:0] tlb__superpage_hits_T_28 = tlb_superpage_entries_2_tag[26:18]; // @[TLB.scala 95:46]
  wire  tlb__superpage_hits_T_30 = tlb__superpage_hits_T_28 == tlb__superpage_hits_T_1; // @[TLB.scala 95:77]
  wire  tlb__superpage_hits_T_32 = tlb_superpage_entries_2_valid_0 & tlb__superpage_hits_T_30; // @[TLB.scala 95:29]
  wire  tlb__superpage_hits_ignore_T_7 = tlb_superpage_entries_2_level < 2'h1; // @[TLB.scala 94:28]
  wire [8:0] tlb__superpage_hits_T_33 = tlb_superpage_entries_2_tag[17:9]; // @[TLB.scala 95:46]
  wire  tlb__superpage_hits_T_35 = tlb__superpage_hits_T_33 == tlb__superpage_hits_T_6; // @[TLB.scala 95:77]
  wire  tlb__superpage_hits_T_36 = tlb__superpage_hits_ignore_T_7 | tlb__superpage_hits_T_35; // @[TLB.scala 95:40]
  wire  tlb__superpage_hits_T_37 = tlb__superpage_hits_T_32 & tlb__superpage_hits_T_36; // @[TLB.scala 95:29]
  wire [8:0] tlb__superpage_hits_T_42 = tlb_superpage_entries_3_tag[26:18]; // @[TLB.scala 95:46]
  wire  tlb__superpage_hits_T_44 = tlb__superpage_hits_T_42 == tlb__superpage_hits_T_1; // @[TLB.scala 95:77]
  wire  tlb__superpage_hits_T_46 = tlb_superpage_entries_3_valid_0 & tlb__superpage_hits_T_44; // @[TLB.scala 95:29]
  wire  tlb__superpage_hits_ignore_T_10 = tlb_superpage_entries_3_level < 2'h1; // @[TLB.scala 94:28]
  wire [8:0] tlb__superpage_hits_T_47 = tlb_superpage_entries_3_tag[17:9]; // @[TLB.scala 95:46]
  wire  tlb__superpage_hits_T_49 = tlb__superpage_hits_T_47 == tlb__superpage_hits_T_6; // @[TLB.scala 95:77]
  wire  tlb__superpage_hits_T_50 = tlb__superpage_hits_ignore_T_10 | tlb__superpage_hits_T_49; // @[TLB.scala 95:40]
  wire  tlb__superpage_hits_T_51 = tlb__superpage_hits_T_46 & tlb__superpage_hits_T_50; // @[TLB.scala 95:29]
  wire [1:0] tlb_hitsVec_idx = tlb_vpn[1:0]; // @[package.scala 143:13]
  wire  tlb__GEN_1 = 2'h1 == tlb_hitsVec_idx ? tlb_sectored_entries_0_valid_1 : tlb_sectored_entries_0_valid_0; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  tlb__GEN_2 = 2'h2 == tlb_hitsVec_idx ? tlb_sectored_entries_0_valid_2 : tlb__GEN_1; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  tlb__GEN_3 = 2'h3 == tlb_hitsVec_idx ? tlb_sectored_entries_0_valid_3 : tlb__GEN_2; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  tlb__hitsVec_T_3 = tlb__GEN_3 & tlb__sector_hits_T_5; // @[TLB.scala 100:18]
  wire  tlb_hitsVec_0 = tlb_vm_enabled & tlb__hitsVec_T_3; // @[TLB.scala 211:44]
  wire  tlb__GEN_5 = 2'h1 == tlb_hitsVec_idx ? tlb_sectored_entries_1_valid_1 : tlb_sectored_entries_1_valid_0; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  tlb__GEN_6 = 2'h2 == tlb_hitsVec_idx ? tlb_sectored_entries_1_valid_2 : tlb__GEN_5; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  tlb__GEN_7 = 2'h3 == tlb_hitsVec_idx ? tlb_sectored_entries_1_valid_3 : tlb__GEN_6; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  tlb__hitsVec_T_7 = tlb__GEN_7 & tlb__sector_hits_T_11; // @[TLB.scala 100:18]
  wire  tlb_hitsVec_1 = tlb_vm_enabled & tlb__hitsVec_T_7; // @[TLB.scala 211:44]
  wire  tlb__GEN_9 = 2'h1 == tlb_hitsVec_idx ? tlb_sectored_entries_2_valid_1 : tlb_sectored_entries_2_valid_0; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  tlb__GEN_10 = 2'h2 == tlb_hitsVec_idx ? tlb_sectored_entries_2_valid_2 : tlb__GEN_9; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  tlb__GEN_11 = 2'h3 == tlb_hitsVec_idx ? tlb_sectored_entries_2_valid_3 : tlb__GEN_10; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  tlb__hitsVec_T_11 = tlb__GEN_11 & tlb__sector_hits_T_17; // @[TLB.scala 100:18]
  wire  tlb_hitsVec_2 = tlb_vm_enabled & tlb__hitsVec_T_11; // @[TLB.scala 211:44]
  wire  tlb__GEN_13 = 2'h1 == tlb_hitsVec_idx ? tlb_sectored_entries_3_valid_1 : tlb_sectored_entries_3_valid_0; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  tlb__GEN_14 = 2'h2 == tlb_hitsVec_idx ? tlb_sectored_entries_3_valid_2 : tlb__GEN_13; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  tlb__GEN_15 = 2'h3 == tlb_hitsVec_idx ? tlb_sectored_entries_3_valid_3 : tlb__GEN_14; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  tlb__hitsVec_T_15 = tlb__GEN_15 & tlb__sector_hits_T_23; // @[TLB.scala 100:18]
  wire  tlb_hitsVec_3 = tlb_vm_enabled & tlb__hitsVec_T_15; // @[TLB.scala 211:44]
  wire  tlb__GEN_17 = 2'h1 == tlb_hitsVec_idx ? tlb_sectored_entries_4_valid_1 : tlb_sectored_entries_4_valid_0; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  tlb__GEN_18 = 2'h2 == tlb_hitsVec_idx ? tlb_sectored_entries_4_valid_2 : tlb__GEN_17; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  tlb__GEN_19 = 2'h3 == tlb_hitsVec_idx ? tlb_sectored_entries_4_valid_3 : tlb__GEN_18; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  tlb__hitsVec_T_19 = tlb__GEN_19 & tlb__sector_hits_T_29; // @[TLB.scala 100:18]
  wire  tlb_hitsVec_4 = tlb_vm_enabled & tlb__hitsVec_T_19; // @[TLB.scala 211:44]
  wire  tlb__GEN_21 = 2'h1 == tlb_hitsVec_idx ? tlb_sectored_entries_5_valid_1 : tlb_sectored_entries_5_valid_0; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  tlb__GEN_22 = 2'h2 == tlb_hitsVec_idx ? tlb_sectored_entries_5_valid_2 : tlb__GEN_21; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  tlb__GEN_23 = 2'h3 == tlb_hitsVec_idx ? tlb_sectored_entries_5_valid_3 : tlb__GEN_22; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  tlb__hitsVec_T_23 = tlb__GEN_23 & tlb__sector_hits_T_35; // @[TLB.scala 100:18]
  wire  tlb_hitsVec_5 = tlb_vm_enabled & tlb__hitsVec_T_23; // @[TLB.scala 211:44]
  wire  tlb__GEN_25 = 2'h1 == tlb_hitsVec_idx ? tlb_sectored_entries_6_valid_1 : tlb_sectored_entries_6_valid_0; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  tlb__GEN_26 = 2'h2 == tlb_hitsVec_idx ? tlb_sectored_entries_6_valid_2 : tlb__GEN_25; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  tlb__GEN_27 = 2'h3 == tlb_hitsVec_idx ? tlb_sectored_entries_6_valid_3 : tlb__GEN_26; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  tlb__hitsVec_T_27 = tlb__GEN_27 & tlb__sector_hits_T_41; // @[TLB.scala 100:18]
  wire  tlb_hitsVec_6 = tlb_vm_enabled & tlb__hitsVec_T_27; // @[TLB.scala 211:44]
  wire  tlb__GEN_29 = 2'h1 == tlb_hitsVec_idx ? tlb_sectored_entries_7_valid_1 : tlb_sectored_entries_7_valid_0; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  tlb__GEN_30 = 2'h2 == tlb_hitsVec_idx ? tlb_sectored_entries_7_valid_2 : tlb__GEN_29; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  tlb__GEN_31 = 2'h3 == tlb_hitsVec_idx ? tlb_sectored_entries_7_valid_3 : tlb__GEN_30; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  tlb__hitsVec_T_31 = tlb__GEN_31 & tlb__sector_hits_T_47; // @[TLB.scala 100:18]
  wire  tlb_hitsVec_7 = tlb_vm_enabled & tlb__hitsVec_T_31; // @[TLB.scala 211:44]
  wire  tlb_hitsVec_8 = tlb_vm_enabled & tlb__superpage_hits_T_9; // @[TLB.scala 211:44]
  wire  tlb_hitsVec_9 = tlb_vm_enabled & tlb__superpage_hits_T_23; // @[TLB.scala 211:44]
  wire  tlb_hitsVec_10 = tlb_vm_enabled & tlb__superpage_hits_T_37; // @[TLB.scala 211:44]
  wire  tlb_hitsVec_11 = tlb_vm_enabled & tlb__superpage_hits_T_51; // @[TLB.scala 211:44]
  wire [8:0] tlb__hitsVec_T_92 = tlb_special_entry_tag[26:18]; // @[TLB.scala 95:46]
  wire  tlb__hitsVec_T_94 = tlb__hitsVec_T_92 == tlb__superpage_hits_T_1; // @[TLB.scala 95:77]
  wire  tlb__hitsVec_T_96 = tlb_special_entry_valid_0 & tlb__hitsVec_T_94; // @[TLB.scala 95:29]
  wire [8:0] tlb__hitsVec_T_97 = tlb_special_entry_tag[17:9]; // @[TLB.scala 95:46]
  wire  tlb__hitsVec_T_99 = tlb__hitsVec_T_97 == tlb__superpage_hits_T_6; // @[TLB.scala 95:77]
  wire  tlb__hitsVec_T_100 = tlb__mpu_ppn_ignore_T | tlb__hitsVec_T_99; // @[TLB.scala 95:40]
  wire  tlb__hitsVec_T_101 = tlb__hitsVec_T_96 & tlb__hitsVec_T_100; // @[TLB.scala 95:29]
  wire [8:0] tlb__hitsVec_T_102 = tlb_special_entry_tag[8:0]; // @[TLB.scala 95:46]
  wire  tlb__hitsVec_T_104 = tlb__hitsVec_T_102 == tlb__superpage_hits_T_11; // @[TLB.scala 95:77]
  wire  tlb__hitsVec_T_105 = tlb__mpu_ppn_ignore_T_1 | tlb__hitsVec_T_104; // @[TLB.scala 95:40]
  wire  tlb__hitsVec_T_106 = tlb__hitsVec_T_101 & tlb__hitsVec_T_105; // @[TLB.scala 95:29]
  wire  tlb_hitsVec_12 = tlb_vm_enabled & tlb__hitsVec_T_106; // @[TLB.scala 211:44]
  wire [5:0] tlb_real_hits_left = {tlb_hitsVec_5,tlb_hitsVec_4,tlb_hitsVec_3,tlb_hitsVec_2,tlb_hitsVec_1,tlb_hitsVec_0}; // @[Cat.scala 29:58]
  wire [12:0] tlb_real_hits = {tlb_hitsVec_12,tlb_hitsVec_11,tlb_hitsVec_10,tlb_hitsVec_9,tlb_hitsVec_8,tlb_hitsVec_7,
    tlb_hitsVec_6,tlb_real_hits_left}; // @[Cat.scala 29:58]
  wire  tlb_hits_right = ~tlb_vm_enabled; // @[TLB.scala 213:18]
  wire [13:0] tlb_hits = {tlb_hits_right,tlb_hitsVec_12,tlb_hitsVec_11,tlb_hitsVec_10,tlb_hitsVec_9,tlb_hitsVec_8,
    tlb_hitsVec_7,tlb_hitsVec_6,tlb_real_hits_left}; // @[Cat.scala 29:58]
  wire [34:0] tlb__GEN_33 = 2'h1 == tlb_hitsVec_idx ? tlb_sectored_entries_0_data_1 : tlb_sectored_entries_0_data_0; // @[]
  wire [34:0] tlb__GEN_34 = 2'h2 == tlb_hitsVec_idx ? tlb_sectored_entries_0_data_2 : tlb__GEN_33; // @[]
  wire [34:0] tlb__GEN_35 = 2'h3 == tlb_hitsVec_idx ? tlb_sectored_entries_0_data_3 : tlb__GEN_34; // @[]
  wire [34:0] tlb__GEN_37 = 2'h1 == tlb_hitsVec_idx ? tlb_sectored_entries_1_data_1 : tlb_sectored_entries_1_data_0; // @[]
  wire [34:0] tlb__GEN_38 = 2'h2 == tlb_hitsVec_idx ? tlb_sectored_entries_1_data_2 : tlb__GEN_37; // @[]
  wire [34:0] tlb__GEN_39 = 2'h3 == tlb_hitsVec_idx ? tlb_sectored_entries_1_data_3 : tlb__GEN_38; // @[]
  wire [34:0] tlb__GEN_41 = 2'h1 == tlb_hitsVec_idx ? tlb_sectored_entries_2_data_1 : tlb_sectored_entries_2_data_0; // @[]
  wire [34:0] tlb__GEN_42 = 2'h2 == tlb_hitsVec_idx ? tlb_sectored_entries_2_data_2 : tlb__GEN_41; // @[]
  wire [34:0] tlb__GEN_43 = 2'h3 == tlb_hitsVec_idx ? tlb_sectored_entries_2_data_3 : tlb__GEN_42; // @[]
  wire [34:0] tlb__GEN_45 = 2'h1 == tlb_hitsVec_idx ? tlb_sectored_entries_3_data_1 : tlb_sectored_entries_3_data_0; // @[]
  wire [34:0] tlb__GEN_46 = 2'h2 == tlb_hitsVec_idx ? tlb_sectored_entries_3_data_2 : tlb__GEN_45; // @[]
  wire [34:0] tlb__GEN_47 = 2'h3 == tlb_hitsVec_idx ? tlb_sectored_entries_3_data_3 : tlb__GEN_46; // @[]
  wire [34:0] tlb__GEN_49 = 2'h1 == tlb_hitsVec_idx ? tlb_sectored_entries_4_data_1 : tlb_sectored_entries_4_data_0; // @[]
  wire [34:0] tlb__GEN_50 = 2'h2 == tlb_hitsVec_idx ? tlb_sectored_entries_4_data_2 : tlb__GEN_49; // @[]
  wire [34:0] tlb__GEN_51 = 2'h3 == tlb_hitsVec_idx ? tlb_sectored_entries_4_data_3 : tlb__GEN_50; // @[]
  wire [34:0] tlb__GEN_53 = 2'h1 == tlb_hitsVec_idx ? tlb_sectored_entries_5_data_1 : tlb_sectored_entries_5_data_0; // @[]
  wire [34:0] tlb__GEN_54 = 2'h2 == tlb_hitsVec_idx ? tlb_sectored_entries_5_data_2 : tlb__GEN_53; // @[]
  wire [34:0] tlb__GEN_55 = 2'h3 == tlb_hitsVec_idx ? tlb_sectored_entries_5_data_3 : tlb__GEN_54; // @[]
  wire [34:0] tlb__GEN_57 = 2'h1 == tlb_hitsVec_idx ? tlb_sectored_entries_6_data_1 : tlb_sectored_entries_6_data_0; // @[]
  wire [34:0] tlb__GEN_58 = 2'h2 == tlb_hitsVec_idx ? tlb_sectored_entries_6_data_2 : tlb__GEN_57; // @[]
  wire [34:0] tlb__GEN_59 = 2'h3 == tlb_hitsVec_idx ? tlb_sectored_entries_6_data_3 : tlb__GEN_58; // @[]
  wire [34:0] tlb__GEN_61 = 2'h1 == tlb_hitsVec_idx ? tlb_sectored_entries_7_data_1 : tlb_sectored_entries_7_data_0; // @[]
  wire [34:0] tlb__GEN_62 = 2'h2 == tlb_hitsVec_idx ? tlb_sectored_entries_7_data_2 : tlb__GEN_61; // @[]
  wire [34:0] tlb__GEN_63 = 2'h3 == tlb_hitsVec_idx ? tlb_sectored_entries_7_data_3 : tlb__GEN_62; // @[]
  wire  tlb__ppn_data_T_149 = tlb_superpage_entries_0_data_0[13]; // @[TLB.scala 86:77]
  wire [1:0] tlb_ppn_right = tlb_ppn_data_barrier_8_io_y_ppn[19:18]; // @[TLB.scala 106:26]
  wire [26:0] tlb__ppn_T_1 = tlb__superpage_hits_ignore_T_1 ? tlb_vpn : 27'h0; // @[TLB.scala 109:28]
  wire [26:0] _GEN_349 = {{7'd0}, tlb_ppn_data_barrier_8_io_y_ppn}; // @[TLB.scala 109:47]
  wire [26:0] tlb__ppn_T_2 = tlb__ppn_T_1 | _GEN_349; // @[TLB.scala 109:47]
  wire [8:0] tlb_ppn_left = tlb__ppn_T_2[17:9]; // @[TLB.scala 109:58]
  wire [26:0] tlb__ppn_T_4 = tlb_vpn | _GEN_349; // @[TLB.scala 109:47]
  wire [8:0] tlb_ppn_left_1 = tlb__ppn_T_4[8:0]; // @[TLB.scala 109:58]
  wire [19:0] tlb__ppn_T_5 = {tlb_ppn_right,tlb_ppn_left,tlb_ppn_left_1}; // @[Cat.scala 29:58]
  wire  tlb__ppn_data_T_165 = tlb_superpage_entries_1_data_0[13]; // @[TLB.scala 86:77]
  wire [1:0] tlb_ppn_right_2 = tlb_ppn_data_barrier_9_io_y_ppn[19:18]; // @[TLB.scala 106:26]
  wire [26:0] tlb__ppn_T_6 = tlb__superpage_hits_ignore_T_4 ? tlb_vpn : 27'h0; // @[TLB.scala 109:28]
  wire [26:0] _GEN_351 = {{7'd0}, tlb_ppn_data_barrier_9_io_y_ppn}; // @[TLB.scala 109:47]
  wire [26:0] tlb__ppn_T_7 = tlb__ppn_T_6 | _GEN_351; // @[TLB.scala 109:47]
  wire [8:0] tlb_ppn_left_2 = tlb__ppn_T_7[17:9]; // @[TLB.scala 109:58]
  wire [26:0] tlb__ppn_T_9 = tlb_vpn | _GEN_351; // @[TLB.scala 109:47]
  wire [8:0] tlb_ppn_left_3 = tlb__ppn_T_9[8:0]; // @[TLB.scala 109:58]
  wire [19:0] tlb__ppn_T_10 = {tlb_ppn_right_2,tlb_ppn_left_2,tlb_ppn_left_3}; // @[Cat.scala 29:58]
  wire  tlb__ppn_data_T_181 = tlb_superpage_entries_2_data_0[13]; // @[TLB.scala 86:77]
  wire [1:0] tlb_ppn_right_4 = tlb_ppn_data_barrier_10_io_y_ppn[19:18]; // @[TLB.scala 106:26]
  wire [26:0] tlb__ppn_T_11 = tlb__superpage_hits_ignore_T_7 ? tlb_vpn : 27'h0; // @[TLB.scala 109:28]
  wire [26:0] _GEN_353 = {{7'd0}, tlb_ppn_data_barrier_10_io_y_ppn}; // @[TLB.scala 109:47]
  wire [26:0] tlb__ppn_T_12 = tlb__ppn_T_11 | _GEN_353; // @[TLB.scala 109:47]
  wire [8:0] tlb_ppn_left_4 = tlb__ppn_T_12[17:9]; // @[TLB.scala 109:58]
  wire [26:0] tlb__ppn_T_14 = tlb_vpn | _GEN_353; // @[TLB.scala 109:47]
  wire [8:0] tlb_ppn_left_5 = tlb__ppn_T_14[8:0]; // @[TLB.scala 109:58]
  wire [19:0] tlb__ppn_T_15 = {tlb_ppn_right_4,tlb_ppn_left_4,tlb_ppn_left_5}; // @[Cat.scala 29:58]
  wire  tlb__ppn_data_T_197 = tlb_superpage_entries_3_data_0[13]; // @[TLB.scala 86:77]
  wire [1:0] tlb_ppn_right_6 = tlb_ppn_data_barrier_11_io_y_ppn[19:18]; // @[TLB.scala 106:26]
  wire [26:0] tlb__ppn_T_16 = tlb__superpage_hits_ignore_T_10 ? tlb_vpn : 27'h0; // @[TLB.scala 109:28]
  wire [26:0] _GEN_355 = {{7'd0}, tlb_ppn_data_barrier_11_io_y_ppn}; // @[TLB.scala 109:47]
  wire [26:0] tlb__ppn_T_17 = tlb__ppn_T_16 | _GEN_355; // @[TLB.scala 109:47]
  wire [8:0] tlb_ppn_left_6 = tlb__ppn_T_17[17:9]; // @[TLB.scala 109:58]
  wire [26:0] tlb__ppn_T_19 = tlb_vpn | _GEN_355; // @[TLB.scala 109:47]
  wire [8:0] tlb_ppn_left_7 = tlb__ppn_T_19[8:0]; // @[TLB.scala 109:58]
  wire [19:0] tlb__ppn_T_20 = {tlb_ppn_right_6,tlb_ppn_left_6,tlb_ppn_left_7}; // @[Cat.scala 29:58]
  wire [1:0] tlb_ppn_right_8 = tlb_ppn_data_barrier_12_io_y_ppn[19:18]; // @[TLB.scala 106:26]
  wire [26:0] _GEN_357 = {{7'd0}, tlb_ppn_data_barrier_12_io_y_ppn}; // @[TLB.scala 109:47]
  wire [26:0] tlb__ppn_T_22 = tlb__mpu_ppn_T_1 | _GEN_357; // @[TLB.scala 109:47]
  wire [8:0] tlb_ppn_left_8 = tlb__ppn_T_22[17:9]; // @[TLB.scala 109:58]
  wire [26:0] tlb__ppn_T_24 = tlb__mpu_ppn_T_3 | _GEN_357; // @[TLB.scala 109:47]
  wire [8:0] tlb_ppn_left_9 = tlb__ppn_T_24[8:0]; // @[TLB.scala 109:58]
  wire [19:0] tlb__ppn_T_25 = {tlb_ppn_right_8,tlb_ppn_left_8,tlb_ppn_left_9}; // @[Cat.scala 29:58]
  wire [19:0] tlb__ppn_T_26 = tlb_vpn[19:0]; // @[TLB.scala 214:77]
  wire [19:0] tlb__ppn_T_27 = tlb_hitsVec_0 ? tlb_ppn_data_barrier_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  wire [19:0] tlb__ppn_T_28 = tlb_hitsVec_1 ? tlb_ppn_data_barrier_1_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  wire [19:0] tlb__ppn_T_29 = tlb_hitsVec_2 ? tlb_ppn_data_barrier_2_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  wire [19:0] tlb__ppn_T_30 = tlb_hitsVec_3 ? tlb_ppn_data_barrier_3_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  wire [19:0] tlb__ppn_T_31 = tlb_hitsVec_4 ? tlb_ppn_data_barrier_4_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  wire [19:0] tlb__ppn_T_32 = tlb_hitsVec_5 ? tlb_ppn_data_barrier_5_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  wire [19:0] tlb__ppn_T_33 = tlb_hitsVec_6 ? tlb_ppn_data_barrier_6_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  wire [19:0] tlb__ppn_T_34 = tlb_hitsVec_7 ? tlb_ppn_data_barrier_7_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  wire [19:0] tlb__ppn_T_35 = tlb_hitsVec_8 ? tlb__ppn_T_5 : 20'h0; // @[Mux.scala 27:72]
  wire [19:0] tlb__ppn_T_36 = tlb_hitsVec_9 ? tlb__ppn_T_10 : 20'h0; // @[Mux.scala 27:72]
  wire [19:0] tlb__ppn_T_37 = tlb_hitsVec_10 ? tlb__ppn_T_15 : 20'h0; // @[Mux.scala 27:72]
  wire [19:0] tlb__ppn_T_38 = tlb_hitsVec_11 ? tlb__ppn_T_20 : 20'h0; // @[Mux.scala 27:72]
  wire [19:0] tlb__ppn_T_39 = tlb_hitsVec_12 ? tlb__ppn_T_25 : 20'h0; // @[Mux.scala 27:72]
  wire [19:0] tlb__ppn_T_40 = tlb_hits_right ? tlb__ppn_T_26 : 20'h0; // @[Mux.scala 27:72]
  wire [19:0] tlb__ppn_T_41 = tlb__ppn_T_27 | tlb__ppn_T_28; // @[Mux.scala 27:72]
  wire [19:0] tlb__ppn_T_42 = tlb__ppn_T_41 | tlb__ppn_T_29; // @[Mux.scala 27:72]
  wire [19:0] tlb__ppn_T_43 = tlb__ppn_T_42 | tlb__ppn_T_30; // @[Mux.scala 27:72]
  wire [19:0] tlb__ppn_T_44 = tlb__ppn_T_43 | tlb__ppn_T_31; // @[Mux.scala 27:72]
  wire [19:0] tlb__ppn_T_45 = tlb__ppn_T_44 | tlb__ppn_T_32; // @[Mux.scala 27:72]
  wire [19:0] tlb__ppn_T_46 = tlb__ppn_T_45 | tlb__ppn_T_33; // @[Mux.scala 27:72]
  wire [19:0] tlb__ppn_T_47 = tlb__ppn_T_46 | tlb__ppn_T_34; // @[Mux.scala 27:72]
  wire [19:0] tlb__ppn_T_48 = tlb__ppn_T_47 | tlb__ppn_T_35; // @[Mux.scala 27:72]
  wire [19:0] tlb__ppn_T_49 = tlb__ppn_T_48 | tlb__ppn_T_36; // @[Mux.scala 27:72]
  wire [19:0] tlb__ppn_T_50 = tlb__ppn_T_49 | tlb__ppn_T_37; // @[Mux.scala 27:72]
  wire [19:0] tlb__ppn_T_51 = tlb__ppn_T_50 | tlb__ppn_T_38; // @[Mux.scala 27:72]
  wire [19:0] tlb__ppn_T_52 = tlb__ppn_T_51 | tlb__ppn_T_39; // @[Mux.scala 27:72]
  wire [19:0] tlb__ppn_T_53 = tlb__ppn_T_52 | tlb__ppn_T_40; // @[Mux.scala 27:72]
  wire  tlb__newEntry_g_T = tlb_io_ptw_resp_bits_pte_g & tlb_io_ptw_resp_bits_pte_v; // @[TLB.scala 223:25]
  wire  tlb__newEntry_sr_T = ~tlb_io_ptw_resp_bits_pte_w; // @[PTW.scala 70:47]
  wire  tlb__newEntry_sr_T_1 = tlb_io_ptw_resp_bits_pte_x & tlb__newEntry_sr_T; // @[PTW.scala 70:44]
  wire  tlb__newEntry_sr_T_2 = tlb_io_ptw_resp_bits_pte_r | tlb__newEntry_sr_T_1; // @[PTW.scala 70:38]
  wire  tlb__newEntry_sr_T_3 = tlb_io_ptw_resp_bits_pte_v & tlb__newEntry_sr_T_2; // @[PTW.scala 70:32]
  wire  tlb__newEntry_sr_T_4 = tlb__newEntry_sr_T_3 & tlb_io_ptw_resp_bits_pte_a; // @[PTW.scala 70:52]
  wire  tlb__newEntry_sr_T_5 = tlb__newEntry_sr_T_4 & tlb_io_ptw_resp_bits_pte_r; // @[PTW.scala 74:35]
  wire  tlb__newEntry_sw_T_5 = tlb__newEntry_sr_T_4 & tlb_io_ptw_resp_bits_pte_w; // @[PTW.scala 75:35]
  wire  tlb__newEntry_sw_T_6 = tlb__newEntry_sw_T_5 & tlb_io_ptw_resp_bits_pte_d; // @[PTW.scala 75:40]
  wire  tlb__newEntry_sx_T_5 = tlb__newEntry_sr_T_4 & tlb_io_ptw_resp_bits_pte_x; // @[PTW.scala 76:35]
  wire  tlb__T = ~tlb_io_ptw_resp_bits_homogeneous; // @[TLB.scala 237:37]
  wire [7:0] tlb_special_entry_data_0_left = {tlb_prot_x,tlb_prot_r,tlb__prot_w_T_31,tlb_prot_al,tlb_prot_al,
    tlb_prot_eff,tlb__cacheable_T_13,1'h0}; // @[TLB.scala 123:24]
  wire [34:0] tlb__special_entry_data_0_T = {tlb_refill_ppn,tlb_io_ptw_resp_bits_pte_u,tlb__newEntry_g_T,
    tlb_io_ptw_resp_bits_ae,tlb__newEntry_sw_T_6,tlb__newEntry_sx_T_5,tlb__newEntry_sr_T_5,tlb_prot_w,
    tlb_special_entry_data_0_left}; // @[TLB.scala 123:24]
  wire  tlb__GEN_64 = tlb_invalidate_refill ? 1'h0 : 1'h1; // @[TLB.scala 240:34 TLB.scala 126:38 TLB.scala 122:16]
  wire  tlb__T_2 = tlb_io_ptw_resp_bits_level < 2'h2; // @[TLB.scala 242:40]
  wire  tlb__T_3 = tlb_r_superpage_repl_addr == 2'h0; // @[TLB.scala 243:82]
  wire  tlb__superpage_entries_0_level_T = tlb_io_ptw_resp_bits_level[0]; // @[package.scala 143:13]
  wire  tlb__GEN_67 = tlb__T_3 ? tlb__GEN_64 : tlb_superpage_entries_0_valid_0; // @[TLB.scala 243:89 TLB.scala 163:30]
  wire  tlb__T_4 = tlb_r_superpage_repl_addr == 2'h1; // @[TLB.scala 243:82]
  wire  tlb__GEN_71 = tlb__T_4 ? tlb__GEN_64 : tlb_superpage_entries_1_valid_0; // @[TLB.scala 243:89 TLB.scala 163:30]
  wire  tlb__T_5 = tlb_r_superpage_repl_addr == 2'h2; // @[TLB.scala 243:82]
  wire  tlb__GEN_75 = tlb__T_5 ? tlb__GEN_64 : tlb_superpage_entries_2_valid_0; // @[TLB.scala 243:89 TLB.scala 163:30]
  wire  tlb__T_6 = tlb_r_superpage_repl_addr == 2'h3; // @[TLB.scala 243:82]
  wire  tlb__GEN_79 = tlb__T_6 ? tlb__GEN_64 : tlb_superpage_entries_3_valid_0; // @[TLB.scala 243:89 TLB.scala 163:30]
  wire [2:0] tlb_waddr = tlb_r_sectored_hit ? tlb_r_sectored_hit_addr : tlb_r_sectored_repl_addr; // @[TLB.scala 248:22]
  wire  tlb__T_7 = tlb_waddr == 3'h0; // @[TLB.scala 249:65]
  wire  tlb__T_8 = ~tlb_r_sectored_hit; // @[TLB.scala 250:15]
  wire  tlb__GEN_81 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_0_valid_0; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  tlb__GEN_82 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_0_valid_1; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  tlb__GEN_83 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_0_valid_2; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  tlb__GEN_84 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_0_valid_3; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire [1:0] tlb_idx = tlb_r_refill_tag[1:0]; // @[package.scala 143:13]
  wire  tlb__GEN_85 = (2'h0 == tlb_idx) | tlb__GEN_81; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  tlb__GEN_86 = (2'h1 == tlb_idx) | tlb__GEN_82; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  tlb__GEN_87 = (2'h2 == tlb_idx) | tlb__GEN_83; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  tlb__GEN_88 = (2'h3 == tlb_idx) | tlb__GEN_84; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire [34:0] tlb__GEN_89 = 2'h0 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_0_data_0; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] tlb__GEN_90 = 2'h1 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_0_data_1; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] tlb__GEN_91 = 2'h2 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_0_data_2; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] tlb__GEN_92 = 2'h3 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_0_data_3; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire  tlb__GEN_93 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_85; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  tlb__GEN_94 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_86; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  tlb__GEN_95 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_87; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  tlb__GEN_96 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_88; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  tlb__GEN_97 = tlb__T_7 ? tlb__GEN_93 : tlb_sectored_entries_0_valid_0; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  tlb__GEN_98 = tlb__T_7 ? tlb__GEN_94 : tlb_sectored_entries_0_valid_1; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  tlb__GEN_99 = tlb__T_7 ? tlb__GEN_95 : tlb_sectored_entries_0_valid_2; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  tlb__GEN_100 = tlb__T_7 ? tlb__GEN_96 : tlb_sectored_entries_0_valid_3; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  tlb__T_9 = tlb_waddr == 3'h1; // @[TLB.scala 249:65]
  wire  tlb__GEN_107 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_1_valid_0; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  tlb__GEN_108 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_1_valid_1; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  tlb__GEN_109 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_1_valid_2; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  tlb__GEN_110 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_1_valid_3; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  tlb__GEN_111 = (2'h0 == tlb_idx) | tlb__GEN_107; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  tlb__GEN_112 = (2'h1 == tlb_idx) | tlb__GEN_108; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  tlb__GEN_113 = (2'h2 == tlb_idx) | tlb__GEN_109; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  tlb__GEN_114 = (2'h3 == tlb_idx) | tlb__GEN_110; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire [34:0] tlb__GEN_115 = 2'h0 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_1_data_0; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] tlb__GEN_116 = 2'h1 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_1_data_1; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] tlb__GEN_117 = 2'h2 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_1_data_2; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] tlb__GEN_118 = 2'h3 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_1_data_3; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire  tlb__GEN_119 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_111; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  tlb__GEN_120 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_112; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  tlb__GEN_121 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_113; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  tlb__GEN_122 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_114; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  tlb__GEN_123 = tlb__T_9 ? tlb__GEN_119 : tlb_sectored_entries_1_valid_0; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  tlb__GEN_124 = tlb__T_9 ? tlb__GEN_120 : tlb_sectored_entries_1_valid_1; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  tlb__GEN_125 = tlb__T_9 ? tlb__GEN_121 : tlb_sectored_entries_1_valid_2; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  tlb__GEN_126 = tlb__T_9 ? tlb__GEN_122 : tlb_sectored_entries_1_valid_3; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  tlb__T_11 = tlb_waddr == 3'h2; // @[TLB.scala 249:65]
  wire  tlb__GEN_133 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_2_valid_0; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  tlb__GEN_134 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_2_valid_1; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  tlb__GEN_135 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_2_valid_2; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  tlb__GEN_136 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_2_valid_3; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  tlb__GEN_137 = (2'h0 == tlb_idx) | tlb__GEN_133; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  tlb__GEN_138 = (2'h1 == tlb_idx) | tlb__GEN_134; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  tlb__GEN_139 = (2'h2 == tlb_idx) | tlb__GEN_135; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  tlb__GEN_140 = (2'h3 == tlb_idx) | tlb__GEN_136; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire [34:0] tlb__GEN_141 = 2'h0 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_2_data_0; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] tlb__GEN_142 = 2'h1 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_2_data_1; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] tlb__GEN_143 = 2'h2 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_2_data_2; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] tlb__GEN_144 = 2'h3 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_2_data_3; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire  tlb__GEN_145 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_137; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  tlb__GEN_146 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_138; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  tlb__GEN_147 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_139; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  tlb__GEN_148 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_140; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  tlb__GEN_149 = tlb__T_11 ? tlb__GEN_145 : tlb_sectored_entries_2_valid_0; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  tlb__GEN_150 = tlb__T_11 ? tlb__GEN_146 : tlb_sectored_entries_2_valid_1; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  tlb__GEN_151 = tlb__T_11 ? tlb__GEN_147 : tlb_sectored_entries_2_valid_2; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  tlb__GEN_152 = tlb__T_11 ? tlb__GEN_148 : tlb_sectored_entries_2_valid_3; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  tlb__T_13 = tlb_waddr == 3'h3; // @[TLB.scala 249:65]
  wire  tlb__GEN_159 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_3_valid_0; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  tlb__GEN_160 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_3_valid_1; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  tlb__GEN_161 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_3_valid_2; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  tlb__GEN_162 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_3_valid_3; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  tlb__GEN_163 = (2'h0 == tlb_idx) | tlb__GEN_159; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  tlb__GEN_164 = (2'h1 == tlb_idx) | tlb__GEN_160; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  tlb__GEN_165 = (2'h2 == tlb_idx) | tlb__GEN_161; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  tlb__GEN_166 = (2'h3 == tlb_idx) | tlb__GEN_162; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire [34:0] tlb__GEN_167 = 2'h0 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_3_data_0; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] tlb__GEN_168 = 2'h1 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_3_data_1; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] tlb__GEN_169 = 2'h2 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_3_data_2; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] tlb__GEN_170 = 2'h3 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_3_data_3; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire  tlb__GEN_171 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_163; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  tlb__GEN_172 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_164; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  tlb__GEN_173 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_165; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  tlb__GEN_174 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_166; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  tlb__GEN_175 = tlb__T_13 ? tlb__GEN_171 : tlb_sectored_entries_3_valid_0; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  tlb__GEN_176 = tlb__T_13 ? tlb__GEN_172 : tlb_sectored_entries_3_valid_1; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  tlb__GEN_177 = tlb__T_13 ? tlb__GEN_173 : tlb_sectored_entries_3_valid_2; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  tlb__GEN_178 = tlb__T_13 ? tlb__GEN_174 : tlb_sectored_entries_3_valid_3; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  tlb__T_15 = tlb_waddr == 3'h4; // @[TLB.scala 249:65]
  wire  tlb__GEN_185 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_4_valid_0; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  tlb__GEN_186 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_4_valid_1; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  tlb__GEN_187 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_4_valid_2; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  tlb__GEN_188 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_4_valid_3; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  tlb__GEN_189 = (2'h0 == tlb_idx) | tlb__GEN_185; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  tlb__GEN_190 = (2'h1 == tlb_idx) | tlb__GEN_186; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  tlb__GEN_191 = (2'h2 == tlb_idx) | tlb__GEN_187; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  tlb__GEN_192 = (2'h3 == tlb_idx) | tlb__GEN_188; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire [34:0] tlb__GEN_193 = 2'h0 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_4_data_0; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] tlb__GEN_194 = 2'h1 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_4_data_1; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] tlb__GEN_195 = 2'h2 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_4_data_2; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] tlb__GEN_196 = 2'h3 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_4_data_3; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire  tlb__GEN_197 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_189; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  tlb__GEN_198 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_190; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  tlb__GEN_199 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_191; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  tlb__GEN_200 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_192; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  tlb__GEN_201 = tlb__T_15 ? tlb__GEN_197 : tlb_sectored_entries_4_valid_0; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  tlb__GEN_202 = tlb__T_15 ? tlb__GEN_198 : tlb_sectored_entries_4_valid_1; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  tlb__GEN_203 = tlb__T_15 ? tlb__GEN_199 : tlb_sectored_entries_4_valid_2; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  tlb__GEN_204 = tlb__T_15 ? tlb__GEN_200 : tlb_sectored_entries_4_valid_3; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  tlb__T_17 = tlb_waddr == 3'h5; // @[TLB.scala 249:65]
  wire  tlb__GEN_211 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_5_valid_0; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  tlb__GEN_212 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_5_valid_1; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  tlb__GEN_213 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_5_valid_2; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  tlb__GEN_214 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_5_valid_3; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  tlb__GEN_215 = (2'h0 == tlb_idx) | tlb__GEN_211; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  tlb__GEN_216 = (2'h1 == tlb_idx) | tlb__GEN_212; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  tlb__GEN_217 = (2'h2 == tlb_idx) | tlb__GEN_213; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  tlb__GEN_218 = (2'h3 == tlb_idx) | tlb__GEN_214; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire [34:0] tlb__GEN_219 = 2'h0 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_5_data_0; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] tlb__GEN_220 = 2'h1 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_5_data_1; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] tlb__GEN_221 = 2'h2 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_5_data_2; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] tlb__GEN_222 = 2'h3 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_5_data_3; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire  tlb__GEN_223 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_215; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  tlb__GEN_224 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_216; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  tlb__GEN_225 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_217; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  tlb__GEN_226 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_218; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  tlb__GEN_227 = tlb__T_17 ? tlb__GEN_223 : tlb_sectored_entries_5_valid_0; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  tlb__GEN_228 = tlb__T_17 ? tlb__GEN_224 : tlb_sectored_entries_5_valid_1; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  tlb__GEN_229 = tlb__T_17 ? tlb__GEN_225 : tlb_sectored_entries_5_valid_2; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  tlb__GEN_230 = tlb__T_17 ? tlb__GEN_226 : tlb_sectored_entries_5_valid_3; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  tlb__T_19 = tlb_waddr == 3'h6; // @[TLB.scala 249:65]
  wire  tlb__GEN_237 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_6_valid_0; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  tlb__GEN_238 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_6_valid_1; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  tlb__GEN_239 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_6_valid_2; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  tlb__GEN_240 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_6_valid_3; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  tlb__GEN_241 = (2'h0 == tlb_idx) | tlb__GEN_237; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  tlb__GEN_242 = (2'h1 == tlb_idx) | tlb__GEN_238; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  tlb__GEN_243 = (2'h2 == tlb_idx) | tlb__GEN_239; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  tlb__GEN_244 = (2'h3 == tlb_idx) | tlb__GEN_240; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire [34:0] tlb__GEN_245 = 2'h0 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_6_data_0; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] tlb__GEN_246 = 2'h1 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_6_data_1; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] tlb__GEN_247 = 2'h2 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_6_data_2; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] tlb__GEN_248 = 2'h3 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_6_data_3; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire  tlb__GEN_249 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_241; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  tlb__GEN_250 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_242; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  tlb__GEN_251 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_243; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  tlb__GEN_252 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_244; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  tlb__GEN_253 = tlb__T_19 ? tlb__GEN_249 : tlb_sectored_entries_6_valid_0; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  tlb__GEN_254 = tlb__T_19 ? tlb__GEN_250 : tlb_sectored_entries_6_valid_1; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  tlb__GEN_255 = tlb__T_19 ? tlb__GEN_251 : tlb_sectored_entries_6_valid_2; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  tlb__GEN_256 = tlb__T_19 ? tlb__GEN_252 : tlb_sectored_entries_6_valid_3; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  tlb__T_21 = tlb_waddr == 3'h7; // @[TLB.scala 249:65]
  wire  tlb__GEN_263 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_7_valid_0; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  tlb__GEN_264 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_7_valid_1; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  tlb__GEN_265 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_7_valid_2; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  tlb__GEN_266 = tlb__T_8 ? 1'h0 : tlb_sectored_entries_7_valid_3; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  tlb__GEN_267 = (2'h0 == tlb_idx) | tlb__GEN_263; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  tlb__GEN_268 = (2'h1 == tlb_idx) | tlb__GEN_264; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  tlb__GEN_269 = (2'h2 == tlb_idx) | tlb__GEN_265; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  tlb__GEN_270 = (2'h3 == tlb_idx) | tlb__GEN_266; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire [34:0] tlb__GEN_271 = 2'h0 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_7_data_0; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] tlb__GEN_272 = 2'h1 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_7_data_1; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] tlb__GEN_273 = 2'h2 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_7_data_2; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] tlb__GEN_274 = 2'h3 == tlb_idx ? tlb__special_entry_data_0_T : tlb_sectored_entries_7_data_3; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire  tlb__GEN_275 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_267; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  tlb__GEN_276 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_268; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  tlb__GEN_277 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_269; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  tlb__GEN_278 = tlb_invalidate_refill ? 1'h0 : tlb__GEN_270; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  tlb__GEN_279 = tlb__T_21 ? tlb__GEN_275 : tlb_sectored_entries_7_valid_0; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  tlb__GEN_280 = tlb__T_21 ? tlb__GEN_276 : tlb_sectored_entries_7_valid_1; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  tlb__GEN_281 = tlb__T_21 ? tlb__GEN_277 : tlb_sectored_entries_7_valid_2; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  tlb__GEN_282 = tlb__T_21 ? tlb__GEN_278 : tlb_sectored_entries_7_valid_3; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  tlb__GEN_291 = tlb__T_2 ? tlb__GEN_67 : tlb_superpage_entries_0_valid_0; // @[TLB.scala 242:54 TLB.scala 163:30]
  wire  tlb__GEN_295 = tlb__T_2 ? tlb__GEN_71 : tlb_superpage_entries_1_valid_0; // @[TLB.scala 242:54 TLB.scala 163:30]
  wire  tlb__GEN_299 = tlb__T_2 ? tlb__GEN_75 : tlb_superpage_entries_2_valid_0; // @[TLB.scala 242:54 TLB.scala 163:30]
  wire  tlb__GEN_303 = tlb__T_2 ? tlb__GEN_79 : tlb_superpage_entries_3_valid_0; // @[TLB.scala 242:54 TLB.scala 163:30]
  wire  tlb__GEN_305 = tlb__T_2 ? tlb_sectored_entries_0_valid_0 : tlb__GEN_97; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  tlb__GEN_306 = tlb__T_2 ? tlb_sectored_entries_0_valid_1 : tlb__GEN_98; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  tlb__GEN_307 = tlb__T_2 ? tlb_sectored_entries_0_valid_2 : tlb__GEN_99; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  tlb__GEN_308 = tlb__T_2 ? tlb_sectored_entries_0_valid_3 : tlb__GEN_100; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  tlb__GEN_315 = tlb__T_2 ? tlb_sectored_entries_1_valid_0 : tlb__GEN_123; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  tlb__GEN_316 = tlb__T_2 ? tlb_sectored_entries_1_valid_1 : tlb__GEN_124; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  tlb__GEN_317 = tlb__T_2 ? tlb_sectored_entries_1_valid_2 : tlb__GEN_125; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  tlb__GEN_318 = tlb__T_2 ? tlb_sectored_entries_1_valid_3 : tlb__GEN_126; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  tlb__GEN_325 = tlb__T_2 ? tlb_sectored_entries_2_valid_0 : tlb__GEN_149; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  tlb__GEN_326 = tlb__T_2 ? tlb_sectored_entries_2_valid_1 : tlb__GEN_150; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  tlb__GEN_327 = tlb__T_2 ? tlb_sectored_entries_2_valid_2 : tlb__GEN_151; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  tlb__GEN_328 = tlb__T_2 ? tlb_sectored_entries_2_valid_3 : tlb__GEN_152; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  tlb__GEN_335 = tlb__T_2 ? tlb_sectored_entries_3_valid_0 : tlb__GEN_175; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  tlb__GEN_336 = tlb__T_2 ? tlb_sectored_entries_3_valid_1 : tlb__GEN_176; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  tlb__GEN_337 = tlb__T_2 ? tlb_sectored_entries_3_valid_2 : tlb__GEN_177; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  tlb__GEN_338 = tlb__T_2 ? tlb_sectored_entries_3_valid_3 : tlb__GEN_178; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  tlb__GEN_345 = tlb__T_2 ? tlb_sectored_entries_4_valid_0 : tlb__GEN_201; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  tlb__GEN_346 = tlb__T_2 ? tlb_sectored_entries_4_valid_1 : tlb__GEN_202; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  tlb__GEN_347 = tlb__T_2 ? tlb_sectored_entries_4_valid_2 : tlb__GEN_203; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  tlb__GEN_348 = tlb__T_2 ? tlb_sectored_entries_4_valid_3 : tlb__GEN_204; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  tlb__GEN_355 = tlb__T_2 ? tlb_sectored_entries_5_valid_0 : tlb__GEN_227; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  tlb__GEN_356 = tlb__T_2 ? tlb_sectored_entries_5_valid_1 : tlb__GEN_228; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  tlb__GEN_357 = tlb__T_2 ? tlb_sectored_entries_5_valid_2 : tlb__GEN_229; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  tlb__GEN_358 = tlb__T_2 ? tlb_sectored_entries_5_valid_3 : tlb__GEN_230; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  tlb__GEN_365 = tlb__T_2 ? tlb_sectored_entries_6_valid_0 : tlb__GEN_253; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  tlb__GEN_366 = tlb__T_2 ? tlb_sectored_entries_6_valid_1 : tlb__GEN_254; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  tlb__GEN_367 = tlb__T_2 ? tlb_sectored_entries_6_valid_2 : tlb__GEN_255; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  tlb__GEN_368 = tlb__T_2 ? tlb_sectored_entries_6_valid_3 : tlb__GEN_256; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  tlb__GEN_375 = tlb__T_2 ? tlb_sectored_entries_7_valid_0 : tlb__GEN_279; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  tlb__GEN_376 = tlb__T_2 ? tlb_sectored_entries_7_valid_1 : tlb__GEN_280; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  tlb__GEN_377 = tlb__T_2 ? tlb_sectored_entries_7_valid_2 : tlb__GEN_281; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  tlb__GEN_378 = tlb__T_2 ? tlb_sectored_entries_7_valid_3 : tlb__GEN_282; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  tlb__GEN_387 = tlb__T ? tlb__GEN_64 : tlb_special_entry_valid_0; // @[TLB.scala 237:68 TLB.scala 164:56]
  wire  tlb__GEN_391 = tlb__T ? tlb_superpage_entries_0_valid_0 : tlb__GEN_291; // @[TLB.scala 237:68 TLB.scala 163:30]
  wire  tlb__GEN_395 = tlb__T ? tlb_superpage_entries_1_valid_0 : tlb__GEN_295; // @[TLB.scala 237:68 TLB.scala 163:30]
  wire  tlb__GEN_399 = tlb__T ? tlb_superpage_entries_2_valid_0 : tlb__GEN_299; // @[TLB.scala 237:68 TLB.scala 163:30]
  wire  tlb__GEN_403 = tlb__T ? tlb_superpage_entries_3_valid_0 : tlb__GEN_303; // @[TLB.scala 237:68 TLB.scala 163:30]
  wire  tlb__GEN_405 = tlb__T ? tlb_sectored_entries_0_valid_0 : tlb__GEN_305; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  tlb__GEN_406 = tlb__T ? tlb_sectored_entries_0_valid_1 : tlb__GEN_306; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  tlb__GEN_407 = tlb__T ? tlb_sectored_entries_0_valid_2 : tlb__GEN_307; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  tlb__GEN_408 = tlb__T ? tlb_sectored_entries_0_valid_3 : tlb__GEN_308; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  tlb__GEN_415 = tlb__T ? tlb_sectored_entries_1_valid_0 : tlb__GEN_315; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  tlb__GEN_416 = tlb__T ? tlb_sectored_entries_1_valid_1 : tlb__GEN_316; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  tlb__GEN_417 = tlb__T ? tlb_sectored_entries_1_valid_2 : tlb__GEN_317; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  tlb__GEN_418 = tlb__T ? tlb_sectored_entries_1_valid_3 : tlb__GEN_318; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  tlb__GEN_425 = tlb__T ? tlb_sectored_entries_2_valid_0 : tlb__GEN_325; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  tlb__GEN_426 = tlb__T ? tlb_sectored_entries_2_valid_1 : tlb__GEN_326; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  tlb__GEN_427 = tlb__T ? tlb_sectored_entries_2_valid_2 : tlb__GEN_327; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  tlb__GEN_428 = tlb__T ? tlb_sectored_entries_2_valid_3 : tlb__GEN_328; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  tlb__GEN_435 = tlb__T ? tlb_sectored_entries_3_valid_0 : tlb__GEN_335; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  tlb__GEN_436 = tlb__T ? tlb_sectored_entries_3_valid_1 : tlb__GEN_336; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  tlb__GEN_437 = tlb__T ? tlb_sectored_entries_3_valid_2 : tlb__GEN_337; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  tlb__GEN_438 = tlb__T ? tlb_sectored_entries_3_valid_3 : tlb__GEN_338; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  tlb__GEN_445 = tlb__T ? tlb_sectored_entries_4_valid_0 : tlb__GEN_345; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  tlb__GEN_446 = tlb__T ? tlb_sectored_entries_4_valid_1 : tlb__GEN_346; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  tlb__GEN_447 = tlb__T ? tlb_sectored_entries_4_valid_2 : tlb__GEN_347; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  tlb__GEN_448 = tlb__T ? tlb_sectored_entries_4_valid_3 : tlb__GEN_348; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  tlb__GEN_455 = tlb__T ? tlb_sectored_entries_5_valid_0 : tlb__GEN_355; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  tlb__GEN_456 = tlb__T ? tlb_sectored_entries_5_valid_1 : tlb__GEN_356; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  tlb__GEN_457 = tlb__T ? tlb_sectored_entries_5_valid_2 : tlb__GEN_357; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  tlb__GEN_458 = tlb__T ? tlb_sectored_entries_5_valid_3 : tlb__GEN_358; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  tlb__GEN_465 = tlb__T ? tlb_sectored_entries_6_valid_0 : tlb__GEN_365; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  tlb__GEN_466 = tlb__T ? tlb_sectored_entries_6_valid_1 : tlb__GEN_366; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  tlb__GEN_467 = tlb__T ? tlb_sectored_entries_6_valid_2 : tlb__GEN_367; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  tlb__GEN_468 = tlb__T ? tlb_sectored_entries_6_valid_3 : tlb__GEN_368; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  tlb__GEN_475 = tlb__T ? tlb_sectored_entries_7_valid_0 : tlb__GEN_375; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  tlb__GEN_476 = tlb__T ? tlb_sectored_entries_7_valid_1 : tlb__GEN_376; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  tlb__GEN_477 = tlb__T ? tlb_sectored_entries_7_valid_2 : tlb__GEN_377; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  tlb__GEN_478 = tlb__T ? tlb_sectored_entries_7_valid_3 : tlb__GEN_378; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  tlb__GEN_487 = tlb_io_ptw_resp_valid ? tlb__GEN_387 : tlb_special_entry_valid_0; // @[TLB.scala 217:20 TLB.scala 164:56]
  wire  tlb__GEN_491 = tlb_io_ptw_resp_valid ? tlb__GEN_391 : tlb_superpage_entries_0_valid_0; // @[TLB.scala 217:20 TLB.scala 163:30]
  wire  tlb__GEN_495 = tlb_io_ptw_resp_valid ? tlb__GEN_395 : tlb_superpage_entries_1_valid_0; // @[TLB.scala 217:20 TLB.scala 163:30]
  wire  tlb__GEN_499 = tlb_io_ptw_resp_valid ? tlb__GEN_399 : tlb_superpage_entries_2_valid_0; // @[TLB.scala 217:20 TLB.scala 163:30]
  wire  tlb__GEN_503 = tlb_io_ptw_resp_valid ? tlb__GEN_403 : tlb_superpage_entries_3_valid_0; // @[TLB.scala 217:20 TLB.scala 163:30]
  wire  tlb__GEN_505 = tlb_io_ptw_resp_valid ? tlb__GEN_405 : tlb_sectored_entries_0_valid_0; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  tlb__GEN_506 = tlb_io_ptw_resp_valid ? tlb__GEN_406 : tlb_sectored_entries_0_valid_1; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  tlb__GEN_507 = tlb_io_ptw_resp_valid ? tlb__GEN_407 : tlb_sectored_entries_0_valid_2; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  tlb__GEN_508 = tlb_io_ptw_resp_valid ? tlb__GEN_408 : tlb_sectored_entries_0_valid_3; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  tlb__GEN_515 = tlb_io_ptw_resp_valid ? tlb__GEN_415 : tlb_sectored_entries_1_valid_0; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  tlb__GEN_516 = tlb_io_ptw_resp_valid ? tlb__GEN_416 : tlb_sectored_entries_1_valid_1; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  tlb__GEN_517 = tlb_io_ptw_resp_valid ? tlb__GEN_417 : tlb_sectored_entries_1_valid_2; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  tlb__GEN_518 = tlb_io_ptw_resp_valid ? tlb__GEN_418 : tlb_sectored_entries_1_valid_3; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  tlb__GEN_525 = tlb_io_ptw_resp_valid ? tlb__GEN_425 : tlb_sectored_entries_2_valid_0; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  tlb__GEN_526 = tlb_io_ptw_resp_valid ? tlb__GEN_426 : tlb_sectored_entries_2_valid_1; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  tlb__GEN_527 = tlb_io_ptw_resp_valid ? tlb__GEN_427 : tlb_sectored_entries_2_valid_2; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  tlb__GEN_528 = tlb_io_ptw_resp_valid ? tlb__GEN_428 : tlb_sectored_entries_2_valid_3; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  tlb__GEN_535 = tlb_io_ptw_resp_valid ? tlb__GEN_435 : tlb_sectored_entries_3_valid_0; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  tlb__GEN_536 = tlb_io_ptw_resp_valid ? tlb__GEN_436 : tlb_sectored_entries_3_valid_1; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  tlb__GEN_537 = tlb_io_ptw_resp_valid ? tlb__GEN_437 : tlb_sectored_entries_3_valid_2; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  tlb__GEN_538 = tlb_io_ptw_resp_valid ? tlb__GEN_438 : tlb_sectored_entries_3_valid_3; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  tlb__GEN_545 = tlb_io_ptw_resp_valid ? tlb__GEN_445 : tlb_sectored_entries_4_valid_0; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  tlb__GEN_546 = tlb_io_ptw_resp_valid ? tlb__GEN_446 : tlb_sectored_entries_4_valid_1; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  tlb__GEN_547 = tlb_io_ptw_resp_valid ? tlb__GEN_447 : tlb_sectored_entries_4_valid_2; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  tlb__GEN_548 = tlb_io_ptw_resp_valid ? tlb__GEN_448 : tlb_sectored_entries_4_valid_3; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  tlb__GEN_555 = tlb_io_ptw_resp_valid ? tlb__GEN_455 : tlb_sectored_entries_5_valid_0; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  tlb__GEN_556 = tlb_io_ptw_resp_valid ? tlb__GEN_456 : tlb_sectored_entries_5_valid_1; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  tlb__GEN_557 = tlb_io_ptw_resp_valid ? tlb__GEN_457 : tlb_sectored_entries_5_valid_2; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  tlb__GEN_558 = tlb_io_ptw_resp_valid ? tlb__GEN_458 : tlb_sectored_entries_5_valid_3; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  tlb__GEN_565 = tlb_io_ptw_resp_valid ? tlb__GEN_465 : tlb_sectored_entries_6_valid_0; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  tlb__GEN_566 = tlb_io_ptw_resp_valid ? tlb__GEN_466 : tlb_sectored_entries_6_valid_1; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  tlb__GEN_567 = tlb_io_ptw_resp_valid ? tlb__GEN_467 : tlb_sectored_entries_6_valid_2; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  tlb__GEN_568 = tlb_io_ptw_resp_valid ? tlb__GEN_468 : tlb_sectored_entries_6_valid_3; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  tlb__GEN_575 = tlb_io_ptw_resp_valid ? tlb__GEN_475 : tlb_sectored_entries_7_valid_0; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  tlb__GEN_576 = tlb_io_ptw_resp_valid ? tlb__GEN_476 : tlb_sectored_entries_7_valid_1; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  tlb__GEN_577 = tlb_io_ptw_resp_valid ? tlb__GEN_477 : tlb_sectored_entries_7_valid_2; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  tlb__GEN_578 = tlb_io_ptw_resp_valid ? tlb__GEN_478 : tlb_sectored_entries_7_valid_3; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire [5:0] tlb_ptw_ae_array_left = {tlb_entries_barrier_5_io_y_ae,tlb_entries_barrier_4_io_y_ae,
    tlb_entries_barrier_3_io_y_ae,tlb_entries_barrier_2_io_y_ae,tlb_entries_barrier_1_io_y_ae,
    tlb_entries_barrier_io_y_ae}; // @[Cat.scala 29:58]
  wire [13:0] tlb_ptw_ae_array = {1'h0,tlb_entries_barrier_12_io_y_ae,tlb_entries_barrier_11_io_y_ae,
    tlb_entries_barrier_10_io_y_ae,tlb_entries_barrier_9_io_y_ae,tlb_entries_barrier_8_io_y_ae,
    tlb_entries_barrier_7_io_y_ae,tlb_entries_barrier_6_io_y_ae,tlb_ptw_ae_array_left}; // @[Cat.scala 29:58]
  wire  tlb__priv_rw_ok_T = ~tlb_priv_s; // @[TLB.scala 261:24]
  wire  tlb__priv_rw_ok_T_1 = tlb__priv_rw_ok_T | tlb_io_ptw_status_sum; // @[TLB.scala 261:32]
  wire [5:0] tlb_priv_rw_ok_left = {tlb_entries_barrier_5_io_y_u,tlb_entries_barrier_4_io_y_u,
    tlb_entries_barrier_3_io_y_u,tlb_entries_barrier_2_io_y_u,tlb_entries_barrier_1_io_y_u,tlb_entries_barrier_io_y_u}; // @[Cat.scala 29:58]
  wire [12:0] tlb__priv_rw_ok_T_2 = {tlb_entries_barrier_12_io_y_u,tlb_entries_barrier_11_io_y_u,
    tlb_entries_barrier_10_io_y_u,tlb_entries_barrier_9_io_y_u,tlb_entries_barrier_8_io_y_u,tlb_entries_barrier_7_io_y_u
    ,tlb_entries_barrier_6_io_y_u,tlb_priv_rw_ok_left}; // @[Cat.scala 29:58]
  wire [12:0] tlb__priv_rw_ok_T_3 = tlb__priv_rw_ok_T_1 ? tlb__priv_rw_ok_T_2 : 13'h0; // @[TLB.scala 261:23]
  wire [12:0] tlb__priv_rw_ok_T_5 = ~tlb__priv_rw_ok_T_2; // @[TLB.scala 261:98]
  wire [12:0] tlb__priv_rw_ok_T_6 = tlb_priv_s ? tlb__priv_rw_ok_T_5 : 13'h0; // @[TLB.scala 261:89]
  wire [12:0] tlb_priv_rw_ok = tlb__priv_rw_ok_T_3 | tlb__priv_rw_ok_T_6; // @[TLB.scala 261:84]
  wire [5:0] tlb_r_array_left = {tlb_entries_barrier_5_io_y_sr,tlb_entries_barrier_4_io_y_sr,
    tlb_entries_barrier_3_io_y_sr,tlb_entries_barrier_2_io_y_sr,tlb_entries_barrier_1_io_y_sr,
    tlb_entries_barrier_io_y_sr}; // @[Cat.scala 29:58]
  wire [12:0] tlb__r_array_T = {tlb_entries_barrier_12_io_y_sr,tlb_entries_barrier_11_io_y_sr,
    tlb_entries_barrier_10_io_y_sr,tlb_entries_barrier_9_io_y_sr,tlb_entries_barrier_8_io_y_sr,
    tlb_entries_barrier_7_io_y_sr,tlb_entries_barrier_6_io_y_sr,tlb_r_array_left}; // @[Cat.scala 29:58]
  wire [5:0] tlb_r_array_left_1 = {tlb_entries_barrier_5_io_y_sx,tlb_entries_barrier_4_io_y_sx,
    tlb_entries_barrier_3_io_y_sx,tlb_entries_barrier_2_io_y_sx,tlb_entries_barrier_1_io_y_sx,
    tlb_entries_barrier_io_y_sx}; // @[Cat.scala 29:58]
  wire [12:0] tlb__r_array_T_1 = {tlb_entries_barrier_12_io_y_sx,tlb_entries_barrier_11_io_y_sx,
    tlb_entries_barrier_10_io_y_sx,tlb_entries_barrier_9_io_y_sx,tlb_entries_barrier_8_io_y_sx,
    tlb_entries_barrier_7_io_y_sx,tlb_entries_barrier_6_io_y_sx,tlb_r_array_left_1}; // @[Cat.scala 29:58]
  wire [12:0] tlb__r_array_T_2 = tlb_io_ptw_status_mxr ? tlb__r_array_T_1 : 13'h0; // @[TLB.scala 263:73]
  wire [12:0] tlb__r_array_T_3 = tlb__r_array_T | tlb__r_array_T_2; // @[TLB.scala 263:68]
  wire [12:0] tlb_r_array_left_2 = tlb_priv_rw_ok & tlb__r_array_T_3; // @[TLB.scala 263:40]
  wire [13:0] tlb_r_array = {1'h1,tlb_r_array_left_2}; // @[Cat.scala 29:58]
  wire [5:0] tlb_w_array_left = {tlb_entries_barrier_5_io_y_sw,tlb_entries_barrier_4_io_y_sw,
    tlb_entries_barrier_3_io_y_sw,tlb_entries_barrier_2_io_y_sw,tlb_entries_barrier_1_io_y_sw,
    tlb_entries_barrier_io_y_sw}; // @[Cat.scala 29:58]
  wire [12:0] tlb__w_array_T = {tlb_entries_barrier_12_io_y_sw,tlb_entries_barrier_11_io_y_sw,
    tlb_entries_barrier_10_io_y_sw,tlb_entries_barrier_9_io_y_sw,tlb_entries_barrier_8_io_y_sw,
    tlb_entries_barrier_7_io_y_sw,tlb_entries_barrier_6_io_y_sw,tlb_w_array_left}; // @[Cat.scala 29:58]
  wire [12:0] tlb_w_array_left_1 = tlb_priv_rw_ok & tlb__w_array_T; // @[TLB.scala 264:40]
  wire [13:0] tlb_w_array = {1'h1,tlb_w_array_left_1}; // @[Cat.scala 29:58]
  wire [1:0] tlb_pr_array_right = tlb_prot_r ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [5:0] tlb_pr_array_left = {tlb_normal_entries_barrier_5_io_y_pr,tlb_normal_entries_barrier_4_io_y_pr,
    tlb_normal_entries_barrier_3_io_y_pr,tlb_normal_entries_barrier_2_io_y_pr,tlb_normal_entries_barrier_1_io_y_pr,
    tlb_normal_entries_barrier_io_y_pr}; // @[Cat.scala 29:58]
  wire [13:0] tlb__pr_array_T_1 = {tlb_pr_array_right,tlb_normal_entries_barrier_11_io_y_pr,
    tlb_normal_entries_barrier_10_io_y_pr,tlb_normal_entries_barrier_9_io_y_pr,tlb_normal_entries_barrier_8_io_y_pr,
    tlb_normal_entries_barrier_7_io_y_pr,tlb_normal_entries_barrier_6_io_y_pr,tlb_pr_array_left}; // @[Cat.scala 29:58]
  wire [13:0] tlb__pr_array_T_2 = ~tlb_ptw_ae_array; // @[TLB.scala 266:89]
  wire [13:0] tlb_pr_array = tlb__pr_array_T_1 & tlb__pr_array_T_2; // @[TLB.scala 266:87]
  wire [1:0] tlb_pw_array_right = tlb_prot_w ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [5:0] tlb_pw_array_left = {tlb_normal_entries_barrier_5_io_y_pw,tlb_normal_entries_barrier_4_io_y_pw,
    tlb_normal_entries_barrier_3_io_y_pw,tlb_normal_entries_barrier_2_io_y_pw,tlb_normal_entries_barrier_1_io_y_pw,
    tlb_normal_entries_barrier_io_y_pw}; // @[Cat.scala 29:58]
  wire [13:0] tlb__pw_array_T_1 = {tlb_pw_array_right,tlb_normal_entries_barrier_11_io_y_pw,
    tlb_normal_entries_barrier_10_io_y_pw,tlb_normal_entries_barrier_9_io_y_pw,tlb_normal_entries_barrier_8_io_y_pw,
    tlb_normal_entries_barrier_7_io_y_pw,tlb_normal_entries_barrier_6_io_y_pw,tlb_pw_array_left}; // @[Cat.scala 29:58]
  wire [13:0] tlb_pw_array = tlb__pw_array_T_1 & tlb__pr_array_T_2; // @[TLB.scala 267:87]
  wire [1:0] tlb_eff_array_right = tlb_prot_eff ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [5:0] tlb_eff_array_left = {tlb_normal_entries_barrier_5_io_y_eff,tlb_normal_entries_barrier_4_io_y_eff,
    tlb_normal_entries_barrier_3_io_y_eff,tlb_normal_entries_barrier_2_io_y_eff,tlb_normal_entries_barrier_1_io_y_eff,
    tlb_normal_entries_barrier_io_y_eff}; // @[Cat.scala 29:58]
  wire [13:0] tlb_eff_array = {tlb_eff_array_right,tlb_normal_entries_barrier_11_io_y_eff,
    tlb_normal_entries_barrier_10_io_y_eff,tlb_normal_entries_barrier_9_io_y_eff,tlb_normal_entries_barrier_8_io_y_eff,
    tlb_normal_entries_barrier_7_io_y_eff,tlb_normal_entries_barrier_6_io_y_eff,tlb_eff_array_left}; // @[Cat.scala 29:58]
  wire [1:0] tlb_c_array_right = tlb__cacheable_T_13 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [5:0] tlb_c_array_left = {tlb_normal_entries_barrier_5_io_y_c,tlb_normal_entries_barrier_4_io_y_c,
    tlb_normal_entries_barrier_3_io_y_c,tlb_normal_entries_barrier_2_io_y_c,tlb_normal_entries_barrier_1_io_y_c,
    tlb_normal_entries_barrier_io_y_c}; // @[Cat.scala 29:58]
  wire [13:0] tlb_c_array = {tlb_c_array_right,tlb_normal_entries_barrier_11_io_y_c,tlb_normal_entries_barrier_10_io_y_c
    ,tlb_normal_entries_barrier_9_io_y_c,tlb_normal_entries_barrier_8_io_y_c,tlb_normal_entries_barrier_7_io_y_c,
    tlb_normal_entries_barrier_6_io_y_c,tlb_c_array_left}; // @[Cat.scala 29:58]
  wire [1:0] tlb_ppp_array_right = tlb__prot_w_T_31 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [5:0] tlb_ppp_array_left = {tlb_normal_entries_barrier_5_io_y_ppp,tlb_normal_entries_barrier_4_io_y_ppp,
    tlb_normal_entries_barrier_3_io_y_ppp,tlb_normal_entries_barrier_2_io_y_ppp,tlb_normal_entries_barrier_1_io_y_ppp,
    tlb_normal_entries_barrier_io_y_ppp}; // @[Cat.scala 29:58]
  wire [13:0] tlb_ppp_array = {tlb_ppp_array_right,tlb_normal_entries_barrier_11_io_y_ppp,
    tlb_normal_entries_barrier_10_io_y_ppp,tlb_normal_entries_barrier_9_io_y_ppp,tlb_normal_entries_barrier_8_io_y_ppp,
    tlb_normal_entries_barrier_7_io_y_ppp,tlb_normal_entries_barrier_6_io_y_ppp,tlb_ppp_array_left}; // @[Cat.scala 29:58]
  wire [1:0] tlb_paa_array_right = tlb_prot_al ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [5:0] tlb_paa_array_left = {tlb_normal_entries_barrier_5_io_y_paa,tlb_normal_entries_barrier_4_io_y_paa,
    tlb_normal_entries_barrier_3_io_y_paa,tlb_normal_entries_barrier_2_io_y_paa,tlb_normal_entries_barrier_1_io_y_paa,
    tlb_normal_entries_barrier_io_y_paa}; // @[Cat.scala 29:58]
  wire [13:0] tlb_paa_array = {tlb_paa_array_right,tlb_normal_entries_barrier_11_io_y_paa,
    tlb_normal_entries_barrier_10_io_y_paa,tlb_normal_entries_barrier_9_io_y_paa,tlb_normal_entries_barrier_8_io_y_paa,
    tlb_normal_entries_barrier_7_io_y_paa,tlb_normal_entries_barrier_6_io_y_paa,tlb_paa_array_left}; // @[Cat.scala 29:58]
  wire [5:0] tlb_pal_array_left = {tlb_normal_entries_barrier_5_io_y_pal,tlb_normal_entries_barrier_4_io_y_pal,
    tlb_normal_entries_barrier_3_io_y_pal,tlb_normal_entries_barrier_2_io_y_pal,tlb_normal_entries_barrier_1_io_y_pal,
    tlb_normal_entries_barrier_io_y_pal}; // @[Cat.scala 29:58]
  wire [13:0] tlb_pal_array = {tlb_paa_array_right,tlb_normal_entries_barrier_11_io_y_pal,
    tlb_normal_entries_barrier_10_io_y_pal,tlb_normal_entries_barrier_9_io_y_pal,tlb_normal_entries_barrier_8_io_y_pal,
    tlb_normal_entries_barrier_7_io_y_pal,tlb_normal_entries_barrier_6_io_y_pal,tlb_pal_array_left}; // @[Cat.scala 29:58]
  wire [13:0] tlb_ppp_array_if_cached = tlb_ppp_array | tlb_c_array; // @[TLB.scala 274:39]
  wire [13:0] tlb_paa_array_if_cached = tlb_paa_array | tlb_c_array; // @[TLB.scala 275:39]
  wire [13:0] tlb_pal_array_if_cached = tlb_pal_array | tlb_c_array; // @[TLB.scala 276:39]
  wire [3:0] tlb__misaligned_T = 4'h1 << tlb_io_req_bits_size; // @[OneHot.scala 58:35]
  wire [3:0] tlb__misaligned_T_2 = tlb__misaligned_T - 4'h1; // @[TLB.scala 279:69]
  wire [39:0] _GEN_391 = {{36'd0}, tlb__misaligned_T_2}; // @[TLB.scala 279:39]
  wire [39:0] tlb__misaligned_T_3 = tlb_io_req_bits_vaddr & _GEN_391; // @[TLB.scala 279:39]
  wire  tlb_misaligned = |tlb__misaligned_T_3; // @[TLB.scala 279:75]
  wire [39:0] tlb_bad_va_maskedVAddr = tlb_io_req_bits_vaddr & 40'hc000000000; // @[TLB.scala 285:43]
  wire  tlb__bad_va_T_1 = tlb_bad_va_maskedVAddr == 40'h0; // @[TLB.scala 286:61]
  wire  tlb__bad_va_T_2 = tlb_bad_va_maskedVAddr == 40'hc000000000; // @[TLB.scala 286:82]
  wire  tlb__bad_va_T_3 = tlb__bad_va_T_1 | tlb__bad_va_T_2; // @[TLB.scala 286:67]
  wire  tlb__bad_va_T_4 = ~tlb__bad_va_T_3; // @[TLB.scala 286:47]
  wire  tlb_bad_va = tlb_vm_enabled & tlb__bad_va_T_4; // @[TLB.scala 280:117]
  wire  tlb__cmd_lrsc_T = tlb_io_req_bits_cmd == 5'h6; // @[package.scala 15:47]
  wire  tlb__cmd_lrsc_T_1 = tlb_io_req_bits_cmd == 5'h7; // @[package.scala 15:47]
  wire  tlb__cmd_lrsc_T_2 = tlb__cmd_lrsc_T | tlb__cmd_lrsc_T_1; // @[package.scala 64:59]
  wire  tlb__cmd_amo_logical_T = tlb_io_req_bits_cmd == 5'h4; // @[package.scala 15:47]
  wire  tlb__cmd_amo_logical_T_1 = tlb_io_req_bits_cmd == 5'h9; // @[package.scala 15:47]
  wire  tlb__cmd_amo_logical_T_2 = tlb_io_req_bits_cmd == 5'ha; // @[package.scala 15:47]
  wire  tlb__cmd_amo_logical_T_3 = tlb_io_req_bits_cmd == 5'hb; // @[package.scala 15:47]
  wire  tlb__cmd_amo_logical_T_4 = tlb__cmd_amo_logical_T | tlb__cmd_amo_logical_T_1; // @[package.scala 64:59]
  wire  tlb__cmd_amo_logical_T_5 = tlb__cmd_amo_logical_T_4 | tlb__cmd_amo_logical_T_2; // @[package.scala 64:59]
  wire  tlb__cmd_amo_logical_T_6 = tlb__cmd_amo_logical_T_5 | tlb__cmd_amo_logical_T_3; // @[package.scala 64:59]
  wire  tlb__cmd_amo_arithmetic_T = tlb_io_req_bits_cmd == 5'h8; // @[package.scala 15:47]
  wire  tlb__cmd_amo_arithmetic_T_1 = tlb_io_req_bits_cmd == 5'hc; // @[package.scala 15:47]
  wire  tlb__cmd_amo_arithmetic_T_2 = tlb_io_req_bits_cmd == 5'hd; // @[package.scala 15:47]
  wire  tlb__cmd_amo_arithmetic_T_3 = tlb_io_req_bits_cmd == 5'he; // @[package.scala 15:47]
  wire  tlb__cmd_amo_arithmetic_T_4 = tlb_io_req_bits_cmd == 5'hf; // @[package.scala 15:47]
  wire  tlb__cmd_amo_arithmetic_T_5 = tlb__cmd_amo_arithmetic_T | tlb__cmd_amo_arithmetic_T_1; // @[package.scala 64:59]
  wire  tlb__cmd_amo_arithmetic_T_6 = tlb__cmd_amo_arithmetic_T_5 | tlb__cmd_amo_arithmetic_T_2; // @[package.scala 64:59]
  wire  tlb__cmd_amo_arithmetic_T_7 = tlb__cmd_amo_arithmetic_T_6 | tlb__cmd_amo_arithmetic_T_3; // @[package.scala 64:59]
  wire  tlb__cmd_amo_arithmetic_T_8 = tlb__cmd_amo_arithmetic_T_7 | tlb__cmd_amo_arithmetic_T_4; // @[package.scala 64:59]
  wire  tlb_cmd_put_partial = tlb_io_req_bits_cmd == 5'h11; // @[TLB.scala 293:41]
  wire  tlb__cmd_read_T = tlb_io_req_bits_cmd == 5'h0; // @[Consts.scala 82:31]
  wire  tlb__cmd_read_T_2 = tlb__cmd_read_T | tlb__cmd_lrsc_T; // @[Consts.scala 82:41]
  wire  tlb__cmd_read_T_4 = tlb__cmd_read_T_2 | tlb__cmd_lrsc_T_1; // @[Consts.scala 82:58]
  wire  tlb__cmd_read_T_21 = tlb__cmd_amo_logical_T_6 | tlb__cmd_amo_arithmetic_T_8; // @[Consts.scala 80:44]
  wire  tlb_cmd_read = tlb__cmd_read_T_4 | tlb__cmd_read_T_21; // @[Consts.scala 82:75]
  wire  tlb__cmd_write_T = tlb_io_req_bits_cmd == 5'h1; // @[Consts.scala 83:32]
  wire  tlb__cmd_write_T_2 = tlb__cmd_write_T | tlb_cmd_put_partial; // @[Consts.scala 83:42]
  wire  tlb__cmd_write_T_4 = tlb__cmd_write_T_2 | tlb__cmd_lrsc_T_1; // @[Consts.scala 83:59]
  wire  tlb_cmd_write = tlb__cmd_write_T_4 | tlb__cmd_read_T_21; // @[Consts.scala 83:76]
  wire  tlb__cmd_write_perms_T = tlb_io_req_bits_cmd == 5'h5; // @[package.scala 15:47]
  wire  tlb__cmd_write_perms_T_1 = tlb_io_req_bits_cmd == 5'h17; // @[package.scala 15:47]
  wire  tlb__cmd_write_perms_T_2 = tlb__cmd_write_perms_T | tlb__cmd_write_perms_T_1; // @[package.scala 64:59]
  wire  tlb_cmd_write_perms = tlb_cmd_write | tlb__cmd_write_perms_T_2; // @[TLB.scala 296:35]
  wire [13:0] tlb__ae_array_T = tlb_misaligned ? tlb_eff_array : 14'h0; // @[TLB.scala 301:8]
  wire [13:0] tlb__ae_array_T_1 = ~tlb_c_array; // @[TLB.scala 302:19]
  wire [13:0] tlb__ae_array_T_2 = tlb__cmd_lrsc_T_2 ? tlb__ae_array_T_1 : 14'h0; // @[TLB.scala 302:8]
  wire [13:0] tlb_ae_array = tlb__ae_array_T | tlb__ae_array_T_2; // @[TLB.scala 301:37]
  wire [13:0] tlb__ae_ld_array_T = ~tlb_pr_array; // @[TLB.scala 303:46]
  wire [13:0] tlb__ae_ld_array_T_1 = tlb_ae_array | tlb__ae_ld_array_T; // @[TLB.scala 303:44]
  wire [13:0] tlb_ae_ld_array = tlb_cmd_read ? tlb__ae_ld_array_T_1 : 14'h0; // @[TLB.scala 303:24]
  wire [13:0] tlb__ae_st_array_T = ~tlb_pw_array; // @[TLB.scala 305:37]
  wire [13:0] tlb__ae_st_array_T_1 = tlb_ae_array | tlb__ae_st_array_T; // @[TLB.scala 305:35]
  wire [13:0] tlb__ae_st_array_T_2 = tlb_cmd_write_perms ? tlb__ae_st_array_T_1 : 14'h0; // @[TLB.scala 305:8]
  wire [13:0] tlb__ae_st_array_T_3 = ~tlb_ppp_array_if_cached; // @[TLB.scala 306:26]
  wire [13:0] tlb__ae_st_array_T_4 = tlb_cmd_put_partial ? tlb__ae_st_array_T_3 : 14'h0; // @[TLB.scala 306:8]
  wire [13:0] tlb__ae_st_array_T_5 = tlb__ae_st_array_T_2 | tlb__ae_st_array_T_4; // @[TLB.scala 305:53]
  wire [13:0] tlb__ae_st_array_T_6 = ~tlb_pal_array_if_cached; // @[TLB.scala 307:26]
  wire [13:0] tlb__ae_st_array_T_7 = tlb__cmd_amo_logical_T_6 ? tlb__ae_st_array_T_6 : 14'h0; // @[TLB.scala 307:8]
  wire [13:0] tlb__ae_st_array_T_8 = tlb__ae_st_array_T_5 | tlb__ae_st_array_T_7; // @[TLB.scala 306:53]
  wire [13:0] tlb__ae_st_array_T_9 = ~tlb_paa_array_if_cached; // @[TLB.scala 308:29]
  wire [13:0] tlb__ae_st_array_T_10 = tlb__cmd_amo_arithmetic_T_8 ? tlb__ae_st_array_T_9 : 14'h0; // @[TLB.scala 308:8]
  wire [13:0] tlb_ae_st_array = tlb__ae_st_array_T_8 | tlb__ae_st_array_T_10; // @[TLB.scala 307:53]
  wire  tlb__ma_ld_array_T = tlb_misaligned & tlb_cmd_read; // @[TLB.scala 314:36]
  wire [13:0] tlb__ma_ld_array_T_1 = ~tlb_eff_array; // @[TLB.scala 314:49]
  wire [13:0] tlb_ma_ld_array = tlb__ma_ld_array_T ? tlb__ma_ld_array_T_1 : 14'h0; // @[TLB.scala 314:24]
  wire  tlb__ma_st_array_T = tlb_misaligned & tlb_cmd_write; // @[TLB.scala 315:36]
  wire [13:0] tlb_ma_st_array = tlb__ma_st_array_T ? tlb__ma_ld_array_T_1 : 14'h0; // @[TLB.scala 315:24]
  wire [13:0] tlb__pf_ld_array_T = tlb_r_array | tlb_ptw_ae_array; // @[TLB.scala 316:45]
  wire [13:0] tlb__pf_ld_array_T_1 = ~tlb__pf_ld_array_T; // @[TLB.scala 316:35]
  wire [13:0] tlb_pf_ld_array = tlb_cmd_read ? tlb__pf_ld_array_T_1 : 14'h0; // @[TLB.scala 316:24]
  wire [13:0] tlb__pf_st_array_T = tlb_w_array | tlb_ptw_ae_array; // @[TLB.scala 317:52]
  wire [13:0] tlb__pf_st_array_T_1 = ~tlb__pf_st_array_T; // @[TLB.scala 317:42]
  wire [13:0] tlb_pf_st_array = tlb_cmd_write_perms ? tlb__pf_st_array_T_1 : 14'h0; // @[TLB.scala 317:24]
  wire  tlb_tlb_hit = |tlb_real_hits; // @[TLB.scala 320:27]
  wire  tlb__tlb_miss_T = ~tlb_bad_va; // @[TLB.scala 321:32]
  wire  tlb__tlb_miss_T_1 = tlb_vm_enabled & tlb__tlb_miss_T; // @[TLB.scala 321:29]
  wire  tlb__tlb_miss_T_2 = ~tlb_tlb_hit; // @[TLB.scala 321:43]
  wire  tlb_tlb_miss = tlb__tlb_miss_T_1 & tlb__tlb_miss_T_2; // @[TLB.scala 321:40]
  reg [6:0] tlb_state_reg; // @[Replacement.scala 158:30]
  reg [2:0] tlb_state_reg_1; // @[Replacement.scala 158:30]
  wire  tlb__T_23 = tlb_io_req_valid & tlb_vm_enabled; // @[TLB.scala 325:22]
  wire  tlb__T_24 = tlb_sector_hits_0 | tlb_sector_hits_1; // @[package.scala 64:59]
  wire  tlb__T_25 = tlb__T_24 | tlb_sector_hits_2; // @[package.scala 64:59]
  wire  tlb__T_26 = tlb__T_25 | tlb_sector_hits_3; // @[package.scala 64:59]
  wire  tlb__T_27 = tlb__T_26 | tlb_sector_hits_4; // @[package.scala 64:59]
  wire  tlb__T_28 = tlb__T_27 | tlb_sector_hits_5; // @[package.scala 64:59]
  wire  tlb__T_29 = tlb__T_28 | tlb_sector_hits_6; // @[package.scala 64:59]
  wire  tlb__T_30 = tlb__T_29 | tlb_sector_hits_7; // @[package.scala 64:59]
  wire [7:0] tlb__T_31 = {tlb_sector_hits_7,tlb_sector_hits_6,tlb_sector_hits_5,tlb_sector_hits_4,tlb_sector_hits_3,
    tlb_sector_hits_2,tlb_sector_hits_1,tlb_sector_hits_0}; // @[Cat.scala 29:58]
  wire [3:0] tlb_hi = tlb__T_31[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] tlb_lo = tlb__T_31[3:0]; // @[OneHot.scala 31:18]
  wire  tlb_right_1 = |tlb_hi; // @[OneHot.scala 32:14]
  wire [3:0] tlb__T_32 = tlb_hi | tlb_lo; // @[OneHot.scala 32:28]
  wire [1:0] tlb_hi_1 = tlb__T_32[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] tlb_lo_1 = tlb__T_32[1:0]; // @[OneHot.scala 31:18]
  wire  tlb_right_2 = |tlb_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] tlb__T_33 = tlb_hi_1 | tlb_lo_1; // @[OneHot.scala 32:28]
  wire  tlb_left_1 = tlb__T_33[1]; // @[CircuitMath.scala 30:8]
  wire [2:0] tlb__T_34 = {tlb_right_1,tlb_right_2,tlb_left_1}; // @[Cat.scala 29:58]
  wire  tlb__state_reg_set_left_older_T = tlb__T_34[2]; // @[Replacement.scala 186:43]
  wire  tlb_state_reg_right_right = ~tlb__state_reg_set_left_older_T; // @[Replacement.scala 186:33]
  wire [2:0] tlb_state_reg_left_subtree_state = tlb_state_reg[5:3]; // @[package.scala 143:13]
  wire [2:0] tlb_state_reg_right_subtree_state = tlb_state_reg[2:0]; // @[Replacement.scala 188:38]
  wire [1:0] tlb__state_reg_T = tlb__T_34[1:0]; // @[package.scala 143:13]
  wire  tlb__state_reg_set_left_older_T_1 = tlb__state_reg_T[1]; // @[Replacement.scala 186:43]
  wire  tlb_state_reg_right_right_1 = ~tlb__state_reg_set_left_older_T_1; // @[Replacement.scala 186:33]
  wire  tlb_state_reg_left_subtree_state_1 = tlb_state_reg_left_subtree_state[1]; // @[package.scala 143:13]
  wire  tlb_state_reg_right_subtree_state_1 = tlb_state_reg_left_subtree_state[0]; // @[Replacement.scala 188:38]
  wire  tlb__state_reg_T_1 = tlb__state_reg_T[0]; // @[package.scala 143:13]
  wire  tlb__state_reg_T_3 = ~tlb__state_reg_T_1; // @[Replacement.scala 208:7]
  wire  tlb_state_reg_right_left = tlb_state_reg_right_right_1 ? tlb_state_reg_left_subtree_state_1 : tlb__state_reg_T_3
    ; // @[Replacement.scala 193:16]
  wire  tlb_state_reg_left = tlb_state_reg_right_right_1 ? tlb__state_reg_T_3 : tlb_state_reg_right_subtree_state_1; // @[Replacement.scala 196:16]
  wire [2:0] tlb__state_reg_T_7 = {tlb_state_reg_right_right_1,tlb_state_reg_right_left,tlb_state_reg_left}; // @[Cat.scala 29:58]
  wire [2:0] tlb_state_reg_right_left_1 = tlb_state_reg_right_right ? tlb_state_reg_left_subtree_state :
    tlb__state_reg_T_7; // @[Replacement.scala 193:16]
  wire  tlb_state_reg_left_subtree_state_2 = tlb_state_reg_right_subtree_state[1]; // @[package.scala 143:13]
  wire  tlb_state_reg_right_subtree_state_2 = tlb_state_reg_right_subtree_state[0]; // @[Replacement.scala 188:38]
  wire  tlb_state_reg_right_left_2 = tlb_state_reg_right_right_1 ? tlb_state_reg_left_subtree_state_2 :
    tlb__state_reg_T_3; // @[Replacement.scala 193:16]
  wire  tlb_state_reg_left_1 = tlb_state_reg_right_right_1 ? tlb__state_reg_T_3 : tlb_state_reg_right_subtree_state_2; // @[Replacement.scala 196:16]
  wire [2:0] tlb__state_reg_T_15 = {tlb_state_reg_right_right_1,tlb_state_reg_right_left_2,tlb_state_reg_left_1}; // @[Cat.scala 29:58]
  wire [2:0] tlb_state_reg_left_2 = tlb_state_reg_right_right ? tlb__state_reg_T_15 : tlb_state_reg_right_subtree_state; // @[Replacement.scala 196:16]
  wire [6:0] tlb__state_reg_T_16 = {tlb_state_reg_right_right,tlb_state_reg_right_left_1,tlb_state_reg_left_2}; // @[Cat.scala 29:58]
  wire  tlb__T_35 = tlb__superpage_hits_T_9 | tlb__superpage_hits_T_23; // @[package.scala 64:59]
  wire  tlb__T_36 = tlb__T_35 | tlb__superpage_hits_T_37; // @[package.scala 64:59]
  wire  tlb__T_37 = tlb__T_36 | tlb__superpage_hits_T_51; // @[package.scala 64:59]
  wire [3:0] tlb__T_38 = {tlb__superpage_hits_T_51,tlb__superpage_hits_T_37,tlb__superpage_hits_T_23,
    tlb__superpage_hits_T_9}; // @[Cat.scala 29:58]
  wire [1:0] tlb_hi_2 = tlb__T_38[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] tlb_lo_2 = tlb__T_38[1:0]; // @[OneHot.scala 31:18]
  wire  tlb_right_4 = |tlb_hi_2; // @[OneHot.scala 32:14]
  wire [1:0] tlb__T_39 = tlb_hi_2 | tlb_lo_2; // @[OneHot.scala 32:28]
  wire  tlb_left_4 = tlb__T_39[1]; // @[CircuitMath.scala 30:8]
  wire [1:0] tlb__T_40 = {tlb_right_4,tlb_left_4}; // @[Cat.scala 29:58]
  wire  tlb__state_reg_1_set_left_older_T = tlb__T_40[1]; // @[Replacement.scala 186:43]
  wire  tlb_state_reg_1_right_right = ~tlb__state_reg_1_set_left_older_T; // @[Replacement.scala 186:33]
  wire  tlb_state_reg_1_left_subtree_state = tlb_state_reg_1[1]; // @[package.scala 143:13]
  wire  tlb_state_reg_1_right_subtree_state = tlb_state_reg_1[0]; // @[Replacement.scala 188:38]
  wire  tlb__state_reg_1_T = tlb__T_40[0]; // @[package.scala 143:13]
  wire  tlb__state_reg_1_T_2 = ~tlb__state_reg_1_T; // @[Replacement.scala 208:7]
  wire  tlb_state_reg_1_right_left = tlb_state_reg_1_right_right ? tlb_state_reg_1_left_subtree_state :
    tlb__state_reg_1_T_2; // @[Replacement.scala 193:16]
  wire  tlb_state_reg_1_left = tlb_state_reg_1_right_right ? tlb__state_reg_1_T_2 : tlb_state_reg_1_right_subtree_state; // @[Replacement.scala 196:16]
  wire [2:0] tlb__state_reg_1_T_6 = {tlb_state_reg_1_right_right,tlb_state_reg_1_right_left,tlb_state_reg_1_left}; // @[Cat.scala 29:58]
  wire [5:0] tlb__multipleHits_T = tlb_real_hits[5:0]; // @[Misc.scala 180:37]
  wire [2:0] tlb__multipleHits_T_1 = tlb__multipleHits_T[2:0]; // @[Misc.scala 180:37]
  wire  tlb__multipleHits_T_2 = tlb__multipleHits_T_1[0]; // @[Misc.scala 180:37]
  wire [1:0] tlb__multipleHits_T_3 = tlb__multipleHits_T_1[2:1]; // @[Misc.scala 181:39]
  wire  tlb__multipleHits_T_4 = tlb__multipleHits_T_3[0]; // @[Misc.scala 180:37]
  wire  tlb__multipleHits_T_5 = tlb__multipleHits_T_3[1]; // @[Misc.scala 181:39]
  wire  tlb_multipleHits_rightOne_1 = tlb__multipleHits_T_4 | tlb__multipleHits_T_5; // @[Misc.scala 182:16]
  wire  tlb__multipleHits_T_7 = tlb__multipleHits_T_4 & tlb__multipleHits_T_5; // @[Misc.scala 182:61]
  wire  tlb_multipleHits_leftOne_2 = tlb__multipleHits_T_2 | tlb_multipleHits_rightOne_1; // @[Misc.scala 182:16]
  wire  tlb__multipleHits_T_9 = tlb__multipleHits_T_2 & tlb_multipleHits_rightOne_1; // @[Misc.scala 182:61]
  wire  tlb_multipleHits_leftTwo = tlb__multipleHits_T_7 | tlb__multipleHits_T_9; // @[Misc.scala 182:49]
  wire [2:0] tlb__multipleHits_T_10 = tlb__multipleHits_T[5:3]; // @[Misc.scala 181:39]
  wire  tlb__multipleHits_T_11 = tlb__multipleHits_T_10[0]; // @[Misc.scala 180:37]
  wire [1:0] tlb__multipleHits_T_12 = tlb__multipleHits_T_10[2:1]; // @[Misc.scala 181:39]
  wire  tlb__multipleHits_T_13 = tlb__multipleHits_T_12[0]; // @[Misc.scala 180:37]
  wire  tlb__multipleHits_T_14 = tlb__multipleHits_T_12[1]; // @[Misc.scala 181:39]
  wire  tlb_multipleHits_rightOne_3 = tlb__multipleHits_T_13 | tlb__multipleHits_T_14; // @[Misc.scala 182:16]
  wire  tlb__multipleHits_T_16 = tlb__multipleHits_T_13 & tlb__multipleHits_T_14; // @[Misc.scala 182:61]
  wire  tlb_multipleHits_rightOne_4 = tlb__multipleHits_T_11 | tlb_multipleHits_rightOne_3; // @[Misc.scala 182:16]
  wire  tlb__multipleHits_T_18 = tlb__multipleHits_T_11 & tlb_multipleHits_rightOne_3; // @[Misc.scala 182:61]
  wire  tlb_multipleHits_rightTwo_2 = tlb__multipleHits_T_16 | tlb__multipleHits_T_18; // @[Misc.scala 182:49]
  wire  tlb_multipleHits_leftOne_5 = tlb_multipleHits_leftOne_2 | tlb_multipleHits_rightOne_4; // @[Misc.scala 182:16]
  wire  tlb__multipleHits_T_19 = tlb_multipleHits_leftTwo | tlb_multipleHits_rightTwo_2; // @[Misc.scala 182:37]
  wire  tlb__multipleHits_T_20 = tlb_multipleHits_leftOne_2 & tlb_multipleHits_rightOne_4; // @[Misc.scala 182:61]
  wire  tlb_multipleHits_leftTwo_1 = tlb__multipleHits_T_19 | tlb__multipleHits_T_20; // @[Misc.scala 182:49]
  wire [6:0] tlb__multipleHits_T_21 = tlb_real_hits[12:6]; // @[Misc.scala 181:39]
  wire [2:0] tlb__multipleHits_T_22 = tlb__multipleHits_T_21[2:0]; // @[Misc.scala 180:37]
  wire  tlb__multipleHits_T_23 = tlb__multipleHits_T_22[0]; // @[Misc.scala 180:37]
  wire [1:0] tlb__multipleHits_T_24 = tlb__multipleHits_T_22[2:1]; // @[Misc.scala 181:39]
  wire  tlb__multipleHits_T_25 = tlb__multipleHits_T_24[0]; // @[Misc.scala 180:37]
  wire  tlb__multipleHits_T_26 = tlb__multipleHits_T_24[1]; // @[Misc.scala 181:39]
  wire  tlb_multipleHits_rightOne_6 = tlb__multipleHits_T_25 | tlb__multipleHits_T_26; // @[Misc.scala 182:16]
  wire  tlb__multipleHits_T_28 = tlb__multipleHits_T_25 & tlb__multipleHits_T_26; // @[Misc.scala 182:61]
  wire  tlb_multipleHits_leftOne_8 = tlb__multipleHits_T_23 | tlb_multipleHits_rightOne_6; // @[Misc.scala 182:16]
  wire  tlb__multipleHits_T_30 = tlb__multipleHits_T_23 & tlb_multipleHits_rightOne_6; // @[Misc.scala 182:61]
  wire  tlb_multipleHits_leftTwo_2 = tlb__multipleHits_T_28 | tlb__multipleHits_T_30; // @[Misc.scala 182:49]
  wire [3:0] tlb__multipleHits_T_31 = tlb__multipleHits_T_21[6:3]; // @[Misc.scala 181:39]
  wire [1:0] tlb__multipleHits_T_32 = tlb__multipleHits_T_31[1:0]; // @[Misc.scala 180:37]
  wire  tlb__multipleHits_T_33 = tlb__multipleHits_T_32[0]; // @[Misc.scala 180:37]
  wire  tlb__multipleHits_T_34 = tlb__multipleHits_T_32[1]; // @[Misc.scala 181:39]
  wire  tlb_multipleHits_leftOne_10 = tlb__multipleHits_T_33 | tlb__multipleHits_T_34; // @[Misc.scala 182:16]
  wire  tlb__multipleHits_T_36 = tlb__multipleHits_T_33 & tlb__multipleHits_T_34; // @[Misc.scala 182:61]
  wire [1:0] tlb__multipleHits_T_37 = tlb__multipleHits_T_31[3:2]; // @[Misc.scala 181:39]
  wire  tlb__multipleHits_T_38 = tlb__multipleHits_T_37[0]; // @[Misc.scala 180:37]
  wire  tlb__multipleHits_T_39 = tlb__multipleHits_T_37[1]; // @[Misc.scala 181:39]
  wire  tlb_multipleHits_rightOne_9 = tlb__multipleHits_T_38 | tlb__multipleHits_T_39; // @[Misc.scala 182:16]
  wire  tlb__multipleHits_T_41 = tlb__multipleHits_T_38 & tlb__multipleHits_T_39; // @[Misc.scala 182:61]
  wire  tlb_multipleHits_rightOne_10 = tlb_multipleHits_leftOne_10 | tlb_multipleHits_rightOne_9; // @[Misc.scala 182:16]
  wire  tlb__multipleHits_T_42 = tlb__multipleHits_T_36 | tlb__multipleHits_T_41; // @[Misc.scala 182:37]
  wire  tlb__multipleHits_T_43 = tlb_multipleHits_leftOne_10 & tlb_multipleHits_rightOne_9; // @[Misc.scala 182:61]
  wire  tlb_multipleHits_rightTwo_5 = tlb__multipleHits_T_42 | tlb__multipleHits_T_43; // @[Misc.scala 182:49]
  wire  tlb_multipleHits_rightOne_11 = tlb_multipleHits_leftOne_8 | tlb_multipleHits_rightOne_10; // @[Misc.scala 182:16]
  wire  tlb__multipleHits_T_44 = tlb_multipleHits_leftTwo_2 | tlb_multipleHits_rightTwo_5; // @[Misc.scala 182:37]
  wire  tlb__multipleHits_T_45 = tlb_multipleHits_leftOne_8 & tlb_multipleHits_rightOne_10; // @[Misc.scala 182:61]
  wire  tlb_multipleHits_rightTwo_6 = tlb__multipleHits_T_44 | tlb__multipleHits_T_45; // @[Misc.scala 182:49]
  wire  tlb__multipleHits_T_47 = tlb_multipleHits_leftTwo_1 | tlb_multipleHits_rightTwo_6; // @[Misc.scala 182:37]
  wire  tlb__multipleHits_T_48 = tlb_multipleHits_leftOne_5 & tlb_multipleHits_rightOne_11; // @[Misc.scala 182:61]
  wire  tlb_multipleHits = tlb__multipleHits_T_47 | tlb__multipleHits_T_48; // @[Misc.scala 182:49]
  wire  tlb__io_resp_pf_ld_T = tlb_bad_va & tlb_cmd_read; // @[TLB.scala 338:28]
  wire [13:0] tlb__io_resp_pf_ld_T_1 = tlb_pf_ld_array & tlb_hits; // @[TLB.scala 338:57]
  wire  tlb__io_resp_pf_ld_T_2 = |tlb__io_resp_pf_ld_T_1; // @[TLB.scala 338:65]
  wire  tlb__io_resp_pf_st_T = tlb_bad_va & tlb_cmd_write_perms; // @[TLB.scala 339:28]
  wire [13:0] tlb__io_resp_pf_st_T_1 = tlb_pf_st_array & tlb_hits; // @[TLB.scala 339:64]
  wire  tlb__io_resp_pf_st_T_2 = |tlb__io_resp_pf_st_T_1; // @[TLB.scala 339:72]
  wire [13:0] tlb__io_resp_ae_ld_T = tlb_ae_ld_array & tlb_hits; // @[TLB.scala 341:33]
  wire [13:0] tlb__io_resp_ae_st_T = tlb_ae_st_array & tlb_hits; // @[TLB.scala 342:33]
  wire [13:0] tlb__io_resp_ma_ld_T = tlb_ma_ld_array & tlb_hits; // @[TLB.scala 344:33]
  wire [13:0] tlb__io_resp_ma_st_T = tlb_ma_st_array & tlb_hits; // @[TLB.scala 345:33]
  wire [13:0] tlb__io_resp_cacheable_T = tlb_c_array & tlb_hits; // @[TLB.scala 347:33]
  wire  tlb__io_resp_miss_T = tlb_io_ptw_resp_valid | tlb_tlb_miss; // @[TLB.scala 350:29]
  wire  tlb__T_41 = tlb_io_req_ready & tlb_io_req_valid; // @[Decoupled.scala 40:37]
  wire  tlb__T_42 = tlb__T_41 & tlb_tlb_miss; // @[TLB.scala 359:25]
  wire  tlb_r_superpage_repl_addr_right = tlb_state_reg_1[2]; // @[Replacement.scala 233:38]
  wire  tlb_r_superpage_repl_addr_left = tlb_r_superpage_repl_addr_right ? tlb_state_reg_1_left_subtree_state :
    tlb_state_reg_1_right_subtree_state; // @[Replacement.scala 240:16]
  wire [1:0] tlb__r_superpage_repl_addr_T_2 = {tlb_r_superpage_repl_addr_right,tlb_r_superpage_repl_addr_left}; // @[Cat.scala 29:58]
  wire [3:0] tlb_r_superpage_repl_addr_valids = {tlb_superpage_entries_3_valid_0,tlb_superpage_entries_2_valid_0,
    tlb_superpage_entries_1_valid_0,tlb_superpage_entries_0_valid_0}; // @[Cat.scala 29:58]
  wire  tlb__r_superpage_repl_addr_T_3 = &tlb_r_superpage_repl_addr_valids; // @[TLB.scala 407:16]
  wire [3:0] tlb__r_superpage_repl_addr_T_4 = ~tlb_r_superpage_repl_addr_valids; // @[TLB.scala 407:43]
  wire  tlb__r_superpage_repl_addr_T_5 = tlb__r_superpage_repl_addr_T_4[0]; // @[OneHot.scala 47:40]
  wire  tlb__r_superpage_repl_addr_T_6 = tlb__r_superpage_repl_addr_T_4[1]; // @[OneHot.scala 47:40]
  wire  tlb__r_superpage_repl_addr_T_7 = tlb__r_superpage_repl_addr_T_4[2]; // @[OneHot.scala 47:40]
  wire [1:0] tlb__r_superpage_repl_addr_T_9 = tlb__r_superpage_repl_addr_T_7 ? 2'h2 : 2'h3; // @[Mux.scala 47:69]
  wire  tlb_r_sectored_repl_addr_right = tlb_state_reg[6]; // @[Replacement.scala 233:38]
  wire  tlb_r_sectored_repl_addr_right_1 = tlb_state_reg_left_subtree_state[2]; // @[Replacement.scala 233:38]
  wire  tlb_r_sectored_repl_addr_left = tlb_r_sectored_repl_addr_right_1 ? tlb_state_reg_left_subtree_state_1 :
    tlb_state_reg_right_subtree_state_1; // @[Replacement.scala 240:16]
  wire [1:0] tlb__r_sectored_repl_addr_T_2 = {tlb_r_sectored_repl_addr_right_1,tlb_r_sectored_repl_addr_left}; // @[Cat.scala 29:58]
  wire  tlb_r_sectored_repl_addr_right_2 = tlb_state_reg_right_subtree_state[2]; // @[Replacement.scala 233:38]
  wire  tlb_r_sectored_repl_addr_left_1 = tlb_r_sectored_repl_addr_right_2 ? tlb_state_reg_left_subtree_state_2 :
    tlb_state_reg_right_subtree_state_2; // @[Replacement.scala 240:16]
  wire [1:0] tlb__r_sectored_repl_addr_T_5 = {tlb_r_sectored_repl_addr_right_2,tlb_r_sectored_repl_addr_left_1}; // @[Cat.scala 29:58]
  wire [1:0] tlb_r_sectored_repl_addr_left_2 = tlb_r_sectored_repl_addr_right ? tlb__r_sectored_repl_addr_T_2 :
    tlb__r_sectored_repl_addr_T_5; // @[Replacement.scala 240:16]
  wire [2:0] tlb__r_sectored_repl_addr_T_6 = {tlb_r_sectored_repl_addr_right,tlb_r_sectored_repl_addr_left_2}; // @[Cat.scala 29:58]
  wire [7:0] tlb_r_sectored_repl_addr_valids = {tlb__sector_hits_T_44,tlb__sector_hits_T_38,tlb__sector_hits_T_32,
    tlb__sector_hits_T_26,tlb__sector_hits_T_20,tlb__sector_hits_T_14,tlb__sector_hits_T_8,tlb__sector_hits_T_2}; // @[Cat.scala 29:58]
  wire  tlb__r_sectored_repl_addr_T_7 = &tlb_r_sectored_repl_addr_valids; // @[TLB.scala 407:16]
  wire [7:0] tlb__r_sectored_repl_addr_T_8 = ~tlb_r_sectored_repl_addr_valids; // @[TLB.scala 407:43]
  wire  tlb__r_sectored_repl_addr_T_9 = tlb__r_sectored_repl_addr_T_8[0]; // @[OneHot.scala 47:40]
  wire  tlb__r_sectored_repl_addr_T_10 = tlb__r_sectored_repl_addr_T_8[1]; // @[OneHot.scala 47:40]
  wire  tlb__r_sectored_repl_addr_T_11 = tlb__r_sectored_repl_addr_T_8[2]; // @[OneHot.scala 47:40]
  wire  tlb__r_sectored_repl_addr_T_12 = tlb__r_sectored_repl_addr_T_8[3]; // @[OneHot.scala 47:40]
  wire  tlb__r_sectored_repl_addr_T_13 = tlb__r_sectored_repl_addr_T_8[4]; // @[OneHot.scala 47:40]
  wire  tlb__r_sectored_repl_addr_T_14 = tlb__r_sectored_repl_addr_T_8[5]; // @[OneHot.scala 47:40]
  wire  tlb__r_sectored_repl_addr_T_15 = tlb__r_sectored_repl_addr_T_8[6]; // @[OneHot.scala 47:40]
  wire [2:0] tlb__r_sectored_repl_addr_T_17 = tlb__r_sectored_repl_addr_T_15 ? 3'h6 : 3'h7; // @[Mux.scala 47:69]
  wire [2:0] tlb__r_sectored_repl_addr_T_18 = tlb__r_sectored_repl_addr_T_14 ? 3'h5 : tlb__r_sectored_repl_addr_T_17; // @[Mux.scala 47:69]
  wire [2:0] tlb__r_sectored_repl_addr_T_19 = tlb__r_sectored_repl_addr_T_13 ? 3'h4 : tlb__r_sectored_repl_addr_T_18; // @[Mux.scala 47:69]
  wire [2:0] tlb__r_sectored_repl_addr_T_20 = tlb__r_sectored_repl_addr_T_12 ? 3'h3 : tlb__r_sectored_repl_addr_T_19; // @[Mux.scala 47:69]
  wire [2:0] tlb__r_sectored_repl_addr_T_21 = tlb__r_sectored_repl_addr_T_11 ? 3'h2 : tlb__r_sectored_repl_addr_T_20; // @[Mux.scala 47:69]
  wire [1:0] tlb__GEN_653 = tlb__T_42 ? 2'h1 : tlb_state; // @[TLB.scala 359:38 TLB.scala 360:13 TLB.scala 169:18]
  wire [1:0] tlb__GEN_659 = tlb_io_sfence_valid ? 2'h0 : tlb__GEN_653; // @[TLB.scala 369:21 TLB.scala 369:29]
  wire [1:0] tlb__state_T = tlb_io_sfence_valid ? 2'h3 : 2'h2; // @[TLB.scala 370:45]
  wire [1:0] tlb__GEN_660 = tlb_io_ptw_req_ready ? tlb__state_T : tlb__GEN_659; // @[TLB.scala 370:31 TLB.scala 370:39]
  wire  tlb__T_44 = tlb_state == 2'h2; // @[TLB.scala 373:17]
  wire  tlb__T_45 = tlb__T_44 & tlb_io_sfence_valid; // @[TLB.scala 373:28]
  wire  tlb__T_46 = ~tlb_io_sfence_bits_rs1; // @[TLB.scala 381:14]
  wire [26:0] tlb__T_47 = tlb_io_sfence_bits_addr[38:12]; // @[TLB.scala 381:58]
  wire  tlb__T_48 = tlb__T_47 == tlb_vpn; // @[TLB.scala 381:72]
  wire  tlb__T_49 = tlb__T_46 | tlb__T_48; // @[TLB.scala 381:34]
  wire  tlb__T_51 = tlb__T_49 | tlb_reset; // @[TLB.scala 381:13]
  wire  tlb__T_52 = ~tlb__T_51; // @[TLB.scala 381:13]
  wire  tlb__GEN_665 = 2'h0 == tlb_hitsVec_idx ? 1'h0 : tlb__GEN_505; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  tlb__GEN_666 = 2'h1 == tlb_hitsVec_idx ? 1'h0 : tlb__GEN_506; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  tlb__GEN_667 = 2'h2 == tlb_hitsVec_idx ? 1'h0 : tlb__GEN_507; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  tlb__GEN_668 = 2'h3 == tlb_hitsVec_idx ? 1'h0 : tlb__GEN_508; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  tlb__GEN_669 = tlb__sector_hits_T_5 ? tlb__GEN_665 : tlb__GEN_505; // @[TLB.scala 131:34]
  wire  tlb__GEN_670 = tlb__sector_hits_T_5 ? tlb__GEN_666 : tlb__GEN_506; // @[TLB.scala 131:34]
  wire  tlb__GEN_671 = tlb__sector_hits_T_5 ? tlb__GEN_667 : tlb__GEN_507; // @[TLB.scala 131:34]
  wire  tlb__GEN_672 = tlb__sector_hits_T_5 ? tlb__GEN_668 : tlb__GEN_508; // @[TLB.scala 131:34]
  wire [8:0] tlb__T_58 = tlb__sector_hits_T_3[26:18]; // @[TLB.scala 135:26]
  wire  tlb__T_59 = tlb__T_58 == 9'h0; // @[TLB.scala 135:61]
  wire  tlb__T_60 = tlb_sectored_entries_0_data_0[0]; // @[TLB.scala 83:39]
  wire  tlb__T_73 = tlb_sectored_entries_0_data_0[13]; // @[TLB.scala 83:39]
  wire  tlb__T_76 = tlb_sectored_entries_0_data_1[0]; // @[TLB.scala 83:39]
  wire  tlb__T_89 = tlb_sectored_entries_0_data_1[13]; // @[TLB.scala 83:39]
  wire  tlb__T_92 = tlb_sectored_entries_0_data_2[0]; // @[TLB.scala 83:39]
  wire  tlb__T_105 = tlb_sectored_entries_0_data_2[13]; // @[TLB.scala 83:39]
  wire  tlb__T_108 = tlb_sectored_entries_0_data_3[0]; // @[TLB.scala 83:39]
  wire  tlb__T_121 = tlb_sectored_entries_0_data_3[13]; // @[TLB.scala 83:39]
  wire  tlb__GEN_673 = tlb__T_60 ? 1'h0 : tlb__GEN_669; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  tlb__GEN_674 = tlb__T_76 ? 1'h0 : tlb__GEN_670; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  tlb__GEN_675 = tlb__T_92 ? 1'h0 : tlb__GEN_671; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  tlb__GEN_676 = tlb__T_108 ? 1'h0 : tlb__GEN_672; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  tlb__T_188 = ~tlb__T_73; // @[TLB.scala 143:13]
  wire  tlb__GEN_681 = tlb__T_188 ? 1'h0 : tlb__GEN_505; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__T_189 = ~tlb__T_89; // @[TLB.scala 143:13]
  wire  tlb__GEN_682 = tlb__T_189 ? 1'h0 : tlb__GEN_506; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__T_190 = ~tlb__T_105; // @[TLB.scala 143:13]
  wire  tlb__GEN_683 = tlb__T_190 ? 1'h0 : tlb__GEN_507; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__T_191 = ~tlb__T_121; // @[TLB.scala 143:13]
  wire  tlb__GEN_684 = tlb__T_191 ? 1'h0 : tlb__GEN_508; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__GEN_685 = tlb_io_sfence_bits_rs2 & tlb__GEN_681; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__GEN_686 = tlb_io_sfence_bits_rs2 & tlb__GEN_682; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__GEN_687 = tlb_io_sfence_bits_rs2 & tlb__GEN_683; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__GEN_688 = tlb_io_sfence_bits_rs2 & tlb__GEN_684; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__GEN_693 = 2'h0 == tlb_hitsVec_idx ? 1'h0 : tlb__GEN_515; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  tlb__GEN_694 = 2'h1 == tlb_hitsVec_idx ? 1'h0 : tlb__GEN_516; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  tlb__GEN_695 = 2'h2 == tlb_hitsVec_idx ? 1'h0 : tlb__GEN_517; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  tlb__GEN_696 = 2'h3 == tlb_hitsVec_idx ? 1'h0 : tlb__GEN_518; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  tlb__GEN_697 = tlb__sector_hits_T_11 ? tlb__GEN_693 : tlb__GEN_515; // @[TLB.scala 131:34]
  wire  tlb__GEN_698 = tlb__sector_hits_T_11 ? tlb__GEN_694 : tlb__GEN_516; // @[TLB.scala 131:34]
  wire  tlb__GEN_699 = tlb__sector_hits_T_11 ? tlb__GEN_695 : tlb__GEN_517; // @[TLB.scala 131:34]
  wire  tlb__GEN_700 = tlb__sector_hits_T_11 ? tlb__GEN_696 : tlb__GEN_518; // @[TLB.scala 131:34]
  wire [8:0] tlb__T_197 = tlb__sector_hits_T_9[26:18]; // @[TLB.scala 135:26]
  wire  tlb__T_198 = tlb__T_197 == 9'h0; // @[TLB.scala 135:61]
  wire  tlb__T_199 = tlb_sectored_entries_1_data_0[0]; // @[TLB.scala 83:39]
  wire  tlb__T_212 = tlb_sectored_entries_1_data_0[13]; // @[TLB.scala 83:39]
  wire  tlb__T_215 = tlb_sectored_entries_1_data_1[0]; // @[TLB.scala 83:39]
  wire  tlb__T_228 = tlb_sectored_entries_1_data_1[13]; // @[TLB.scala 83:39]
  wire  tlb__T_231 = tlb_sectored_entries_1_data_2[0]; // @[TLB.scala 83:39]
  wire  tlb__T_244 = tlb_sectored_entries_1_data_2[13]; // @[TLB.scala 83:39]
  wire  tlb__T_247 = tlb_sectored_entries_1_data_3[0]; // @[TLB.scala 83:39]
  wire  tlb__T_260 = tlb_sectored_entries_1_data_3[13]; // @[TLB.scala 83:39]
  wire  tlb__GEN_701 = tlb__T_199 ? 1'h0 : tlb__GEN_697; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  tlb__GEN_702 = tlb__T_215 ? 1'h0 : tlb__GEN_698; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  tlb__GEN_703 = tlb__T_231 ? 1'h0 : tlb__GEN_699; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  tlb__GEN_704 = tlb__T_247 ? 1'h0 : tlb__GEN_700; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  tlb__T_327 = ~tlb__T_212; // @[TLB.scala 143:13]
  wire  tlb__GEN_709 = tlb__T_327 ? 1'h0 : tlb__GEN_515; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__T_328 = ~tlb__T_228; // @[TLB.scala 143:13]
  wire  tlb__GEN_710 = tlb__T_328 ? 1'h0 : tlb__GEN_516; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__T_329 = ~tlb__T_244; // @[TLB.scala 143:13]
  wire  tlb__GEN_711 = tlb__T_329 ? 1'h0 : tlb__GEN_517; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__T_330 = ~tlb__T_260; // @[TLB.scala 143:13]
  wire  tlb__GEN_712 = tlb__T_330 ? 1'h0 : tlb__GEN_518; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__GEN_713 = tlb_io_sfence_bits_rs2 & tlb__GEN_709; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__GEN_714 = tlb_io_sfence_bits_rs2 & tlb__GEN_710; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__GEN_715 = tlb_io_sfence_bits_rs2 & tlb__GEN_711; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__GEN_716 = tlb_io_sfence_bits_rs2 & tlb__GEN_712; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__GEN_721 = 2'h0 == tlb_hitsVec_idx ? 1'h0 : tlb__GEN_525; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  tlb__GEN_722 = 2'h1 == tlb_hitsVec_idx ? 1'h0 : tlb__GEN_526; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  tlb__GEN_723 = 2'h2 == tlb_hitsVec_idx ? 1'h0 : tlb__GEN_527; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  tlb__GEN_724 = 2'h3 == tlb_hitsVec_idx ? 1'h0 : tlb__GEN_528; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  tlb__GEN_725 = tlb__sector_hits_T_17 ? tlb__GEN_721 : tlb__GEN_525; // @[TLB.scala 131:34]
  wire  tlb__GEN_726 = tlb__sector_hits_T_17 ? tlb__GEN_722 : tlb__GEN_526; // @[TLB.scala 131:34]
  wire  tlb__GEN_727 = tlb__sector_hits_T_17 ? tlb__GEN_723 : tlb__GEN_527; // @[TLB.scala 131:34]
  wire  tlb__GEN_728 = tlb__sector_hits_T_17 ? tlb__GEN_724 : tlb__GEN_528; // @[TLB.scala 131:34]
  wire [8:0] tlb__T_336 = tlb__sector_hits_T_15[26:18]; // @[TLB.scala 135:26]
  wire  tlb__T_337 = tlb__T_336 == 9'h0; // @[TLB.scala 135:61]
  wire  tlb__T_338 = tlb_sectored_entries_2_data_0[0]; // @[TLB.scala 83:39]
  wire  tlb__T_351 = tlb_sectored_entries_2_data_0[13]; // @[TLB.scala 83:39]
  wire  tlb__T_354 = tlb_sectored_entries_2_data_1[0]; // @[TLB.scala 83:39]
  wire  tlb__T_367 = tlb_sectored_entries_2_data_1[13]; // @[TLB.scala 83:39]
  wire  tlb__T_370 = tlb_sectored_entries_2_data_2[0]; // @[TLB.scala 83:39]
  wire  tlb__T_383 = tlb_sectored_entries_2_data_2[13]; // @[TLB.scala 83:39]
  wire  tlb__T_386 = tlb_sectored_entries_2_data_3[0]; // @[TLB.scala 83:39]
  wire  tlb__T_399 = tlb_sectored_entries_2_data_3[13]; // @[TLB.scala 83:39]
  wire  tlb__GEN_729 = tlb__T_338 ? 1'h0 : tlb__GEN_725; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  tlb__GEN_730 = tlb__T_354 ? 1'h0 : tlb__GEN_726; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  tlb__GEN_731 = tlb__T_370 ? 1'h0 : tlb__GEN_727; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  tlb__GEN_732 = tlb__T_386 ? 1'h0 : tlb__GEN_728; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  tlb__T_466 = ~tlb__T_351; // @[TLB.scala 143:13]
  wire  tlb__GEN_737 = tlb__T_466 ? 1'h0 : tlb__GEN_525; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__T_467 = ~tlb__T_367; // @[TLB.scala 143:13]
  wire  tlb__GEN_738 = tlb__T_467 ? 1'h0 : tlb__GEN_526; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__T_468 = ~tlb__T_383; // @[TLB.scala 143:13]
  wire  tlb__GEN_739 = tlb__T_468 ? 1'h0 : tlb__GEN_527; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__T_469 = ~tlb__T_399; // @[TLB.scala 143:13]
  wire  tlb__GEN_740 = tlb__T_469 ? 1'h0 : tlb__GEN_528; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__GEN_741 = tlb_io_sfence_bits_rs2 & tlb__GEN_737; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__GEN_742 = tlb_io_sfence_bits_rs2 & tlb__GEN_738; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__GEN_743 = tlb_io_sfence_bits_rs2 & tlb__GEN_739; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__GEN_744 = tlb_io_sfence_bits_rs2 & tlb__GEN_740; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__GEN_749 = 2'h0 == tlb_hitsVec_idx ? 1'h0 : tlb__GEN_535; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  tlb__GEN_750 = 2'h1 == tlb_hitsVec_idx ? 1'h0 : tlb__GEN_536; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  tlb__GEN_751 = 2'h2 == tlb_hitsVec_idx ? 1'h0 : tlb__GEN_537; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  tlb__GEN_752 = 2'h3 == tlb_hitsVec_idx ? 1'h0 : tlb__GEN_538; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  tlb__GEN_753 = tlb__sector_hits_T_23 ? tlb__GEN_749 : tlb__GEN_535; // @[TLB.scala 131:34]
  wire  tlb__GEN_754 = tlb__sector_hits_T_23 ? tlb__GEN_750 : tlb__GEN_536; // @[TLB.scala 131:34]
  wire  tlb__GEN_755 = tlb__sector_hits_T_23 ? tlb__GEN_751 : tlb__GEN_537; // @[TLB.scala 131:34]
  wire  tlb__GEN_756 = tlb__sector_hits_T_23 ? tlb__GEN_752 : tlb__GEN_538; // @[TLB.scala 131:34]
  wire [8:0] tlb__T_475 = tlb__sector_hits_T_21[26:18]; // @[TLB.scala 135:26]
  wire  tlb__T_476 = tlb__T_475 == 9'h0; // @[TLB.scala 135:61]
  wire  tlb__T_477 = tlb_sectored_entries_3_data_0[0]; // @[TLB.scala 83:39]
  wire  tlb__T_490 = tlb_sectored_entries_3_data_0[13]; // @[TLB.scala 83:39]
  wire  tlb__T_493 = tlb_sectored_entries_3_data_1[0]; // @[TLB.scala 83:39]
  wire  tlb__T_506 = tlb_sectored_entries_3_data_1[13]; // @[TLB.scala 83:39]
  wire  tlb__T_509 = tlb_sectored_entries_3_data_2[0]; // @[TLB.scala 83:39]
  wire  tlb__T_522 = tlb_sectored_entries_3_data_2[13]; // @[TLB.scala 83:39]
  wire  tlb__T_525 = tlb_sectored_entries_3_data_3[0]; // @[TLB.scala 83:39]
  wire  tlb__T_538 = tlb_sectored_entries_3_data_3[13]; // @[TLB.scala 83:39]
  wire  tlb__GEN_757 = tlb__T_477 ? 1'h0 : tlb__GEN_753; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  tlb__GEN_758 = tlb__T_493 ? 1'h0 : tlb__GEN_754; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  tlb__GEN_759 = tlb__T_509 ? 1'h0 : tlb__GEN_755; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  tlb__GEN_760 = tlb__T_525 ? 1'h0 : tlb__GEN_756; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  tlb__T_605 = ~tlb__T_490; // @[TLB.scala 143:13]
  wire  tlb__GEN_765 = tlb__T_605 ? 1'h0 : tlb__GEN_535; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__T_606 = ~tlb__T_506; // @[TLB.scala 143:13]
  wire  tlb__GEN_766 = tlb__T_606 ? 1'h0 : tlb__GEN_536; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__T_607 = ~tlb__T_522; // @[TLB.scala 143:13]
  wire  tlb__GEN_767 = tlb__T_607 ? 1'h0 : tlb__GEN_537; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__T_608 = ~tlb__T_538; // @[TLB.scala 143:13]
  wire  tlb__GEN_768 = tlb__T_608 ? 1'h0 : tlb__GEN_538; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__GEN_769 = tlb_io_sfence_bits_rs2 & tlb__GEN_765; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__GEN_770 = tlb_io_sfence_bits_rs2 & tlb__GEN_766; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__GEN_771 = tlb_io_sfence_bits_rs2 & tlb__GEN_767; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__GEN_772 = tlb_io_sfence_bits_rs2 & tlb__GEN_768; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__GEN_777 = 2'h0 == tlb_hitsVec_idx ? 1'h0 : tlb__GEN_545; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  tlb__GEN_778 = 2'h1 == tlb_hitsVec_idx ? 1'h0 : tlb__GEN_546; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  tlb__GEN_779 = 2'h2 == tlb_hitsVec_idx ? 1'h0 : tlb__GEN_547; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  tlb__GEN_780 = 2'h3 == tlb_hitsVec_idx ? 1'h0 : tlb__GEN_548; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  tlb__GEN_781 = tlb__sector_hits_T_29 ? tlb__GEN_777 : tlb__GEN_545; // @[TLB.scala 131:34]
  wire  tlb__GEN_782 = tlb__sector_hits_T_29 ? tlb__GEN_778 : tlb__GEN_546; // @[TLB.scala 131:34]
  wire  tlb__GEN_783 = tlb__sector_hits_T_29 ? tlb__GEN_779 : tlb__GEN_547; // @[TLB.scala 131:34]
  wire  tlb__GEN_784 = tlb__sector_hits_T_29 ? tlb__GEN_780 : tlb__GEN_548; // @[TLB.scala 131:34]
  wire [8:0] tlb__T_614 = tlb__sector_hits_T_27[26:18]; // @[TLB.scala 135:26]
  wire  tlb__T_615 = tlb__T_614 == 9'h0; // @[TLB.scala 135:61]
  wire  tlb__T_616 = tlb_sectored_entries_4_data_0[0]; // @[TLB.scala 83:39]
  wire  tlb__T_629 = tlb_sectored_entries_4_data_0[13]; // @[TLB.scala 83:39]
  wire  tlb__T_632 = tlb_sectored_entries_4_data_1[0]; // @[TLB.scala 83:39]
  wire  tlb__T_645 = tlb_sectored_entries_4_data_1[13]; // @[TLB.scala 83:39]
  wire  tlb__T_648 = tlb_sectored_entries_4_data_2[0]; // @[TLB.scala 83:39]
  wire  tlb__T_661 = tlb_sectored_entries_4_data_2[13]; // @[TLB.scala 83:39]
  wire  tlb__T_664 = tlb_sectored_entries_4_data_3[0]; // @[TLB.scala 83:39]
  wire  tlb__T_677 = tlb_sectored_entries_4_data_3[13]; // @[TLB.scala 83:39]
  wire  tlb__GEN_785 = tlb__T_616 ? 1'h0 : tlb__GEN_781; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  tlb__GEN_786 = tlb__T_632 ? 1'h0 : tlb__GEN_782; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  tlb__GEN_787 = tlb__T_648 ? 1'h0 : tlb__GEN_783; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  tlb__GEN_788 = tlb__T_664 ? 1'h0 : tlb__GEN_784; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  tlb__T_744 = ~tlb__T_629; // @[TLB.scala 143:13]
  wire  tlb__GEN_793 = tlb__T_744 ? 1'h0 : tlb__GEN_545; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__T_745 = ~tlb__T_645; // @[TLB.scala 143:13]
  wire  tlb__GEN_794 = tlb__T_745 ? 1'h0 : tlb__GEN_546; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__T_746 = ~tlb__T_661; // @[TLB.scala 143:13]
  wire  tlb__GEN_795 = tlb__T_746 ? 1'h0 : tlb__GEN_547; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__T_747 = ~tlb__T_677; // @[TLB.scala 143:13]
  wire  tlb__GEN_796 = tlb__T_747 ? 1'h0 : tlb__GEN_548; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__GEN_797 = tlb_io_sfence_bits_rs2 & tlb__GEN_793; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__GEN_798 = tlb_io_sfence_bits_rs2 & tlb__GEN_794; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__GEN_799 = tlb_io_sfence_bits_rs2 & tlb__GEN_795; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__GEN_800 = tlb_io_sfence_bits_rs2 & tlb__GEN_796; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__GEN_805 = 2'h0 == tlb_hitsVec_idx ? 1'h0 : tlb__GEN_555; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  tlb__GEN_806 = 2'h1 == tlb_hitsVec_idx ? 1'h0 : tlb__GEN_556; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  tlb__GEN_807 = 2'h2 == tlb_hitsVec_idx ? 1'h0 : tlb__GEN_557; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  tlb__GEN_808 = 2'h3 == tlb_hitsVec_idx ? 1'h0 : tlb__GEN_558; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  tlb__GEN_809 = tlb__sector_hits_T_35 ? tlb__GEN_805 : tlb__GEN_555; // @[TLB.scala 131:34]
  wire  tlb__GEN_810 = tlb__sector_hits_T_35 ? tlb__GEN_806 : tlb__GEN_556; // @[TLB.scala 131:34]
  wire  tlb__GEN_811 = tlb__sector_hits_T_35 ? tlb__GEN_807 : tlb__GEN_557; // @[TLB.scala 131:34]
  wire  tlb__GEN_812 = tlb__sector_hits_T_35 ? tlb__GEN_808 : tlb__GEN_558; // @[TLB.scala 131:34]
  wire [8:0] tlb__T_753 = tlb__sector_hits_T_33[26:18]; // @[TLB.scala 135:26]
  wire  tlb__T_754 = tlb__T_753 == 9'h0; // @[TLB.scala 135:61]
  wire  tlb__T_755 = tlb_sectored_entries_5_data_0[0]; // @[TLB.scala 83:39]
  wire  tlb__T_768 = tlb_sectored_entries_5_data_0[13]; // @[TLB.scala 83:39]
  wire  tlb__T_771 = tlb_sectored_entries_5_data_1[0]; // @[TLB.scala 83:39]
  wire  tlb__T_784 = tlb_sectored_entries_5_data_1[13]; // @[TLB.scala 83:39]
  wire  tlb__T_787 = tlb_sectored_entries_5_data_2[0]; // @[TLB.scala 83:39]
  wire  tlb__T_800 = tlb_sectored_entries_5_data_2[13]; // @[TLB.scala 83:39]
  wire  tlb__T_803 = tlb_sectored_entries_5_data_3[0]; // @[TLB.scala 83:39]
  wire  tlb__T_816 = tlb_sectored_entries_5_data_3[13]; // @[TLB.scala 83:39]
  wire  tlb__GEN_813 = tlb__T_755 ? 1'h0 : tlb__GEN_809; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  tlb__GEN_814 = tlb__T_771 ? 1'h0 : tlb__GEN_810; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  tlb__GEN_815 = tlb__T_787 ? 1'h0 : tlb__GEN_811; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  tlb__GEN_816 = tlb__T_803 ? 1'h0 : tlb__GEN_812; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  tlb__T_883 = ~tlb__T_768; // @[TLB.scala 143:13]
  wire  tlb__GEN_821 = tlb__T_883 ? 1'h0 : tlb__GEN_555; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__T_884 = ~tlb__T_784; // @[TLB.scala 143:13]
  wire  tlb__GEN_822 = tlb__T_884 ? 1'h0 : tlb__GEN_556; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__T_885 = ~tlb__T_800; // @[TLB.scala 143:13]
  wire  tlb__GEN_823 = tlb__T_885 ? 1'h0 : tlb__GEN_557; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__T_886 = ~tlb__T_816; // @[TLB.scala 143:13]
  wire  tlb__GEN_824 = tlb__T_886 ? 1'h0 : tlb__GEN_558; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__GEN_825 = tlb_io_sfence_bits_rs2 & tlb__GEN_821; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__GEN_826 = tlb_io_sfence_bits_rs2 & tlb__GEN_822; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__GEN_827 = tlb_io_sfence_bits_rs2 & tlb__GEN_823; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__GEN_828 = tlb_io_sfence_bits_rs2 & tlb__GEN_824; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__GEN_833 = 2'h0 == tlb_hitsVec_idx ? 1'h0 : tlb__GEN_565; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  tlb__GEN_834 = 2'h1 == tlb_hitsVec_idx ? 1'h0 : tlb__GEN_566; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  tlb__GEN_835 = 2'h2 == tlb_hitsVec_idx ? 1'h0 : tlb__GEN_567; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  tlb__GEN_836 = 2'h3 == tlb_hitsVec_idx ? 1'h0 : tlb__GEN_568; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  tlb__GEN_837 = tlb__sector_hits_T_41 ? tlb__GEN_833 : tlb__GEN_565; // @[TLB.scala 131:34]
  wire  tlb__GEN_838 = tlb__sector_hits_T_41 ? tlb__GEN_834 : tlb__GEN_566; // @[TLB.scala 131:34]
  wire  tlb__GEN_839 = tlb__sector_hits_T_41 ? tlb__GEN_835 : tlb__GEN_567; // @[TLB.scala 131:34]
  wire  tlb__GEN_840 = tlb__sector_hits_T_41 ? tlb__GEN_836 : tlb__GEN_568; // @[TLB.scala 131:34]
  wire [8:0] tlb__T_892 = tlb__sector_hits_T_39[26:18]; // @[TLB.scala 135:26]
  wire  tlb__T_893 = tlb__T_892 == 9'h0; // @[TLB.scala 135:61]
  wire  tlb__T_894 = tlb_sectored_entries_6_data_0[0]; // @[TLB.scala 83:39]
  wire  tlb__T_907 = tlb_sectored_entries_6_data_0[13]; // @[TLB.scala 83:39]
  wire  tlb__T_910 = tlb_sectored_entries_6_data_1[0]; // @[TLB.scala 83:39]
  wire  tlb__T_923 = tlb_sectored_entries_6_data_1[13]; // @[TLB.scala 83:39]
  wire  tlb__T_926 = tlb_sectored_entries_6_data_2[0]; // @[TLB.scala 83:39]
  wire  tlb__T_939 = tlb_sectored_entries_6_data_2[13]; // @[TLB.scala 83:39]
  wire  tlb__T_942 = tlb_sectored_entries_6_data_3[0]; // @[TLB.scala 83:39]
  wire  tlb__T_955 = tlb_sectored_entries_6_data_3[13]; // @[TLB.scala 83:39]
  wire  tlb__GEN_841 = tlb__T_894 ? 1'h0 : tlb__GEN_837; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  tlb__GEN_842 = tlb__T_910 ? 1'h0 : tlb__GEN_838; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  tlb__GEN_843 = tlb__T_926 ? 1'h0 : tlb__GEN_839; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  tlb__GEN_844 = tlb__T_942 ? 1'h0 : tlb__GEN_840; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  tlb__T_1022 = ~tlb__T_907; // @[TLB.scala 143:13]
  wire  tlb__GEN_849 = tlb__T_1022 ? 1'h0 : tlb__GEN_565; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__T_1023 = ~tlb__T_923; // @[TLB.scala 143:13]
  wire  tlb__GEN_850 = tlb__T_1023 ? 1'h0 : tlb__GEN_566; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__T_1024 = ~tlb__T_939; // @[TLB.scala 143:13]
  wire  tlb__GEN_851 = tlb__T_1024 ? 1'h0 : tlb__GEN_567; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__T_1025 = ~tlb__T_955; // @[TLB.scala 143:13]
  wire  tlb__GEN_852 = tlb__T_1025 ? 1'h0 : tlb__GEN_568; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__GEN_853 = tlb_io_sfence_bits_rs2 & tlb__GEN_849; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__GEN_854 = tlb_io_sfence_bits_rs2 & tlb__GEN_850; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__GEN_855 = tlb_io_sfence_bits_rs2 & tlb__GEN_851; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__GEN_856 = tlb_io_sfence_bits_rs2 & tlb__GEN_852; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__GEN_861 = 2'h0 == tlb_hitsVec_idx ? 1'h0 : tlb__GEN_575; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  tlb__GEN_862 = 2'h1 == tlb_hitsVec_idx ? 1'h0 : tlb__GEN_576; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  tlb__GEN_863 = 2'h2 == tlb_hitsVec_idx ? 1'h0 : tlb__GEN_577; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  tlb__GEN_864 = 2'h3 == tlb_hitsVec_idx ? 1'h0 : tlb__GEN_578; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  tlb__GEN_865 = tlb__sector_hits_T_47 ? tlb__GEN_861 : tlb__GEN_575; // @[TLB.scala 131:34]
  wire  tlb__GEN_866 = tlb__sector_hits_T_47 ? tlb__GEN_862 : tlb__GEN_576; // @[TLB.scala 131:34]
  wire  tlb__GEN_867 = tlb__sector_hits_T_47 ? tlb__GEN_863 : tlb__GEN_577; // @[TLB.scala 131:34]
  wire  tlb__GEN_868 = tlb__sector_hits_T_47 ? tlb__GEN_864 : tlb__GEN_578; // @[TLB.scala 131:34]
  wire [8:0] tlb__T_1031 = tlb__sector_hits_T_45[26:18]; // @[TLB.scala 135:26]
  wire  tlb__T_1032 = tlb__T_1031 == 9'h0; // @[TLB.scala 135:61]
  wire  tlb__T_1033 = tlb_sectored_entries_7_data_0[0]; // @[TLB.scala 83:39]
  wire  tlb__T_1046 = tlb_sectored_entries_7_data_0[13]; // @[TLB.scala 83:39]
  wire  tlb__T_1049 = tlb_sectored_entries_7_data_1[0]; // @[TLB.scala 83:39]
  wire  tlb__T_1062 = tlb_sectored_entries_7_data_1[13]; // @[TLB.scala 83:39]
  wire  tlb__T_1065 = tlb_sectored_entries_7_data_2[0]; // @[TLB.scala 83:39]
  wire  tlb__T_1078 = tlb_sectored_entries_7_data_2[13]; // @[TLB.scala 83:39]
  wire  tlb__T_1081 = tlb_sectored_entries_7_data_3[0]; // @[TLB.scala 83:39]
  wire  tlb__T_1094 = tlb_sectored_entries_7_data_3[13]; // @[TLB.scala 83:39]
  wire  tlb__GEN_869 = tlb__T_1033 ? 1'h0 : tlb__GEN_865; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  tlb__GEN_870 = tlb__T_1049 ? 1'h0 : tlb__GEN_866; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  tlb__GEN_871 = tlb__T_1065 ? 1'h0 : tlb__GEN_867; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  tlb__GEN_872 = tlb__T_1081 ? 1'h0 : tlb__GEN_868; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  tlb__T_1161 = ~tlb__T_1046; // @[TLB.scala 143:13]
  wire  tlb__GEN_877 = tlb__T_1161 ? 1'h0 : tlb__GEN_575; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__T_1162 = ~tlb__T_1062; // @[TLB.scala 143:13]
  wire  tlb__GEN_878 = tlb__T_1162 ? 1'h0 : tlb__GEN_576; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__T_1163 = ~tlb__T_1078; // @[TLB.scala 143:13]
  wire  tlb__GEN_879 = tlb__T_1163 ? 1'h0 : tlb__GEN_577; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__T_1164 = ~tlb__T_1094; // @[TLB.scala 143:13]
  wire  tlb__GEN_880 = tlb__T_1164 ? 1'h0 : tlb__GEN_578; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__GEN_881 = tlb_io_sfence_bits_rs2 & tlb__GEN_877; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__GEN_882 = tlb_io_sfence_bits_rs2 & tlb__GEN_878; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__GEN_883 = tlb_io_sfence_bits_rs2 & tlb__GEN_879; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__GEN_884 = tlb_io_sfence_bits_rs2 & tlb__GEN_880; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__T_1196 = ~tlb__ppn_data_T_149; // @[TLB.scala 143:13]
  wire  tlb__GEN_890 = tlb__T_1196 ? 1'h0 : tlb__GEN_491; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__GEN_891 = tlb_io_sfence_bits_rs2 & tlb__GEN_890; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__T_1228 = ~tlb__ppn_data_T_165; // @[TLB.scala 143:13]
  wire  tlb__GEN_894 = tlb__T_1228 ? 1'h0 : tlb__GEN_495; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__GEN_895 = tlb_io_sfence_bits_rs2 & tlb__GEN_894; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__T_1260 = ~tlb__ppn_data_T_181; // @[TLB.scala 143:13]
  wire  tlb__GEN_898 = tlb__T_1260 ? 1'h0 : tlb__GEN_499; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__GEN_899 = tlb_io_sfence_bits_rs2 & tlb__GEN_898; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__T_1292 = ~tlb__ppn_data_T_197; // @[TLB.scala 143:13]
  wire  tlb__GEN_902 = tlb__T_1292 ? 1'h0 : tlb__GEN_503; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__GEN_903 = tlb_io_sfence_bits_rs2 & tlb__GEN_902; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__T_1324 = ~tlb__mpu_ppn_data_T_13; // @[TLB.scala 143:13]
  wire  tlb__GEN_906 = tlb__T_1324 ? 1'h0 : tlb__GEN_487; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  tlb__GEN_907 = tlb_io_sfence_bits_rs2 & tlb__GEN_906; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  tlb__T_1326 = tlb_multipleHits | tlb_reset; // @[TLB.scala 388:24]
  wire [1:0] pma_checker_io_req_bits_size;
  wire [19:0] pma_checker_mpu_ppn_data_barrier_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_mpu_ppn_data_barrier_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_mpu_ppn_data_barrier_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_mpu_ppn_data_barrier_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_mpu_ppn_data_barrier_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_mpu_ppn_data_barrier_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_mpu_ppn_data_barrier_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_mpu_ppn_data_barrier_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_mpu_ppn_data_barrier_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_mpu_ppn_data_barrier_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_mpu_ppn_data_barrier_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_mpu_ppn_data_barrier_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_mpu_ppn_data_barrier_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_mpu_ppn_data_barrier_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_mpu_ppn_data_barrier_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_mpu_ppn_data_barrier_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_mpu_ppn_data_barrier_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_mpu_ppn_data_barrier_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_mpu_ppn_data_barrier_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_mpu_ppn_data_barrier_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_mpu_ppn_data_barrier_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_mpu_ppn_data_barrier_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_mpu_ppn_data_barrier_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_mpu_ppn_data_barrier_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_mpu_ppn_data_barrier_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_mpu_ppn_data_barrier_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_mpu_ppn_data_barrier_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_mpu_ppn_data_barrier_io_y_c; // @[package.scala 236:25]
  wire [1:0] pma_checker_pmp_io_prv; // @[TLB.scala 190:19]
  wire  pma_checker_pmp_io_pmp_0_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pma_checker_pmp_io_pmp_0_cfg_a; // @[TLB.scala 190:19]
  wire  pma_checker_pmp_io_pmp_0_cfg_x; // @[TLB.scala 190:19]
  wire  pma_checker_pmp_io_pmp_0_cfg_w; // @[TLB.scala 190:19]
  wire  pma_checker_pmp_io_pmp_0_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pma_checker_pmp_io_pmp_0_addr; // @[TLB.scala 190:19]
  wire [31:0] pma_checker_pmp_io_pmp_0_mask; // @[TLB.scala 190:19]
  wire  pma_checker_pmp_io_pmp_1_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pma_checker_pmp_io_pmp_1_cfg_a; // @[TLB.scala 190:19]
  wire  pma_checker_pmp_io_pmp_1_cfg_x; // @[TLB.scala 190:19]
  wire  pma_checker_pmp_io_pmp_1_cfg_w; // @[TLB.scala 190:19]
  wire  pma_checker_pmp_io_pmp_1_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pma_checker_pmp_io_pmp_1_addr; // @[TLB.scala 190:19]
  wire [31:0] pma_checker_pmp_io_pmp_1_mask; // @[TLB.scala 190:19]
  wire  pma_checker_pmp_io_pmp_2_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pma_checker_pmp_io_pmp_2_cfg_a; // @[TLB.scala 190:19]
  wire  pma_checker_pmp_io_pmp_2_cfg_x; // @[TLB.scala 190:19]
  wire  pma_checker_pmp_io_pmp_2_cfg_w; // @[TLB.scala 190:19]
  wire  pma_checker_pmp_io_pmp_2_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pma_checker_pmp_io_pmp_2_addr; // @[TLB.scala 190:19]
  wire [31:0] pma_checker_pmp_io_pmp_2_mask; // @[TLB.scala 190:19]
  wire  pma_checker_pmp_io_pmp_3_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pma_checker_pmp_io_pmp_3_cfg_a; // @[TLB.scala 190:19]
  wire  pma_checker_pmp_io_pmp_3_cfg_x; // @[TLB.scala 190:19]
  wire  pma_checker_pmp_io_pmp_3_cfg_w; // @[TLB.scala 190:19]
  wire  pma_checker_pmp_io_pmp_3_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pma_checker_pmp_io_pmp_3_addr; // @[TLB.scala 190:19]
  wire [31:0] pma_checker_pmp_io_pmp_3_mask; // @[TLB.scala 190:19]
  wire  pma_checker_pmp_io_pmp_4_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pma_checker_pmp_io_pmp_4_cfg_a; // @[TLB.scala 190:19]
  wire  pma_checker_pmp_io_pmp_4_cfg_x; // @[TLB.scala 190:19]
  wire  pma_checker_pmp_io_pmp_4_cfg_w; // @[TLB.scala 190:19]
  wire  pma_checker_pmp_io_pmp_4_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pma_checker_pmp_io_pmp_4_addr; // @[TLB.scala 190:19]
  wire [31:0] pma_checker_pmp_io_pmp_4_mask; // @[TLB.scala 190:19]
  wire  pma_checker_pmp_io_pmp_5_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pma_checker_pmp_io_pmp_5_cfg_a; // @[TLB.scala 190:19]
  wire  pma_checker_pmp_io_pmp_5_cfg_x; // @[TLB.scala 190:19]
  wire  pma_checker_pmp_io_pmp_5_cfg_w; // @[TLB.scala 190:19]
  wire  pma_checker_pmp_io_pmp_5_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pma_checker_pmp_io_pmp_5_addr; // @[TLB.scala 190:19]
  wire [31:0] pma_checker_pmp_io_pmp_5_mask; // @[TLB.scala 190:19]
  wire  pma_checker_pmp_io_pmp_6_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pma_checker_pmp_io_pmp_6_cfg_a; // @[TLB.scala 190:19]
  wire  pma_checker_pmp_io_pmp_6_cfg_x; // @[TLB.scala 190:19]
  wire  pma_checker_pmp_io_pmp_6_cfg_w; // @[TLB.scala 190:19]
  wire  pma_checker_pmp_io_pmp_6_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pma_checker_pmp_io_pmp_6_addr; // @[TLB.scala 190:19]
  wire [31:0] pma_checker_pmp_io_pmp_6_mask; // @[TLB.scala 190:19]
  wire  pma_checker_pmp_io_pmp_7_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pma_checker_pmp_io_pmp_7_cfg_a; // @[TLB.scala 190:19]
  wire  pma_checker_pmp_io_pmp_7_cfg_x; // @[TLB.scala 190:19]
  wire  pma_checker_pmp_io_pmp_7_cfg_w; // @[TLB.scala 190:19]
  wire  pma_checker_pmp_io_pmp_7_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pma_checker_pmp_io_pmp_7_addr; // @[TLB.scala 190:19]
  wire [31:0] pma_checker_pmp_io_pmp_7_mask; // @[TLB.scala 190:19]
  wire [31:0] pma_checker_pmp_io_addr; // @[TLB.scala 190:19]
  wire [1:0] pma_checker_pmp_io_size; // @[TLB.scala 190:19]
  wire  pma_checker_pmp_io_r; // @[TLB.scala 190:19]
  wire  pma_checker_pmp_io_w; // @[TLB.scala 190:19]
  wire  pma_checker_pmp_io_x; // @[TLB.scala 190:19]
  wire [19:0] pma_checker_ppn_data_barrier_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_ppn_data_barrier_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_ppn_data_barrier_1_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_1_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_1_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_1_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_1_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_1_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_1_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_1_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_1_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_1_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_1_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_1_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_1_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_1_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_ppn_data_barrier_1_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_1_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_1_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_1_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_1_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_1_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_1_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_1_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_1_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_1_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_1_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_1_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_1_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_1_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_ppn_data_barrier_2_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_2_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_2_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_2_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_2_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_2_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_2_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_2_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_2_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_2_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_2_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_2_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_2_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_2_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_ppn_data_barrier_2_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_2_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_2_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_2_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_2_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_2_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_2_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_2_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_2_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_2_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_2_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_2_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_2_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_2_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_ppn_data_barrier_3_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_3_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_3_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_3_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_3_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_3_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_3_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_3_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_3_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_3_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_3_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_3_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_3_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_3_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_ppn_data_barrier_3_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_3_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_3_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_3_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_3_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_3_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_3_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_3_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_3_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_3_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_3_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_3_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_3_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_3_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_ppn_data_barrier_4_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_4_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_4_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_4_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_4_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_4_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_4_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_4_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_4_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_4_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_4_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_4_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_4_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_4_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_ppn_data_barrier_4_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_4_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_4_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_4_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_4_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_4_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_4_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_4_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_4_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_4_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_4_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_4_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_4_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_4_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_ppn_data_barrier_5_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_5_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_5_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_5_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_5_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_5_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_5_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_5_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_5_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_5_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_5_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_5_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_5_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_5_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_ppn_data_barrier_5_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_5_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_5_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_5_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_5_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_5_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_5_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_5_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_5_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_5_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_5_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_5_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_5_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_5_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_ppn_data_barrier_6_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_6_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_6_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_6_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_6_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_6_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_6_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_6_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_6_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_6_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_6_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_6_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_6_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_6_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_ppn_data_barrier_6_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_6_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_6_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_6_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_6_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_6_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_6_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_6_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_6_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_6_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_6_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_6_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_6_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_6_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_ppn_data_barrier_7_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_7_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_7_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_7_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_7_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_7_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_7_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_7_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_7_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_7_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_7_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_7_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_7_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_7_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_ppn_data_barrier_7_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_7_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_7_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_7_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_7_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_7_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_7_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_7_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_7_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_7_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_7_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_7_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_7_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_7_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_ppn_data_barrier_8_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_8_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_8_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_8_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_8_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_8_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_8_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_8_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_8_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_8_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_8_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_8_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_8_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_8_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_ppn_data_barrier_8_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_8_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_8_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_8_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_8_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_8_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_8_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_8_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_8_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_8_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_8_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_8_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_8_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_8_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_ppn_data_barrier_9_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_9_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_9_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_9_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_9_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_9_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_9_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_9_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_9_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_9_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_9_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_9_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_9_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_9_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_ppn_data_barrier_9_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_9_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_9_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_9_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_9_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_9_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_9_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_9_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_9_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_9_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_9_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_9_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_9_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_9_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_ppn_data_barrier_10_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_10_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_10_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_10_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_10_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_10_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_10_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_10_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_10_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_10_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_10_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_10_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_10_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_10_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_ppn_data_barrier_10_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_10_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_10_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_10_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_10_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_10_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_10_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_10_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_10_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_10_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_10_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_10_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_10_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_10_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_ppn_data_barrier_11_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_11_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_11_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_11_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_11_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_11_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_11_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_11_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_11_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_11_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_11_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_11_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_11_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_11_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_ppn_data_barrier_11_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_11_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_11_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_11_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_11_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_11_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_11_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_11_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_11_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_11_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_11_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_11_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_11_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_11_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_ppn_data_barrier_12_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_12_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_12_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_12_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_12_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_12_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_12_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_12_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_12_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_12_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_12_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_12_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_12_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_12_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_ppn_data_barrier_12_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_12_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_12_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_12_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_12_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_12_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_12_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_12_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_12_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_12_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_12_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_12_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_12_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_ppn_data_barrier_12_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_entries_barrier_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_entries_barrier_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_entries_barrier_1_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_1_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_1_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_1_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_1_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_1_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_1_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_1_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_1_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_1_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_1_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_1_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_1_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_1_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_entries_barrier_1_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_1_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_1_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_1_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_1_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_1_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_1_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_1_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_1_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_1_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_1_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_1_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_1_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_1_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_entries_barrier_2_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_2_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_2_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_2_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_2_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_2_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_2_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_2_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_2_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_2_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_2_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_2_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_2_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_2_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_entries_barrier_2_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_2_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_2_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_2_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_2_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_2_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_2_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_2_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_2_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_2_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_2_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_2_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_2_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_2_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_entries_barrier_3_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_3_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_3_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_3_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_3_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_3_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_3_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_3_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_3_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_3_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_3_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_3_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_3_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_3_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_entries_barrier_3_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_3_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_3_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_3_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_3_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_3_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_3_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_3_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_3_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_3_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_3_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_3_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_3_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_3_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_entries_barrier_4_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_4_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_4_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_4_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_4_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_4_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_4_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_4_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_4_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_4_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_4_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_4_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_4_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_4_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_entries_barrier_4_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_4_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_4_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_4_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_4_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_4_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_4_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_4_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_4_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_4_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_4_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_4_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_4_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_4_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_entries_barrier_5_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_5_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_5_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_5_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_5_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_5_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_5_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_5_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_5_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_5_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_5_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_5_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_5_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_5_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_entries_barrier_5_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_5_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_5_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_5_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_5_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_5_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_5_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_5_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_5_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_5_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_5_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_5_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_5_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_5_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_entries_barrier_6_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_6_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_6_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_6_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_6_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_6_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_6_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_6_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_6_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_6_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_6_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_6_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_6_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_6_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_entries_barrier_6_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_6_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_6_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_6_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_6_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_6_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_6_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_6_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_6_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_6_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_6_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_6_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_6_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_6_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_entries_barrier_7_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_7_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_7_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_7_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_7_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_7_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_7_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_7_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_7_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_7_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_7_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_7_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_7_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_7_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_entries_barrier_7_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_7_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_7_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_7_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_7_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_7_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_7_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_7_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_7_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_7_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_7_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_7_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_7_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_7_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_entries_barrier_8_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_8_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_8_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_8_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_8_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_8_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_8_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_8_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_8_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_8_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_8_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_8_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_8_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_8_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_entries_barrier_8_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_8_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_8_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_8_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_8_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_8_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_8_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_8_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_8_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_8_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_8_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_8_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_8_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_8_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_entries_barrier_9_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_9_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_9_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_9_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_9_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_9_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_9_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_9_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_9_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_9_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_9_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_9_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_9_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_9_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_entries_barrier_9_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_9_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_9_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_9_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_9_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_9_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_9_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_9_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_9_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_9_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_9_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_9_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_9_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_9_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_entries_barrier_10_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_10_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_10_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_10_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_10_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_10_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_10_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_10_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_10_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_10_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_10_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_10_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_10_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_10_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_entries_barrier_10_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_10_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_10_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_10_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_10_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_10_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_10_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_10_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_10_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_10_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_10_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_10_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_10_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_10_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_entries_barrier_11_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_11_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_11_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_11_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_11_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_11_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_11_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_11_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_11_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_11_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_11_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_11_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_11_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_11_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_entries_barrier_11_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_11_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_11_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_11_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_11_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_11_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_11_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_11_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_11_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_11_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_11_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_11_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_11_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_11_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_entries_barrier_12_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_12_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_12_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_12_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_12_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_12_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_12_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_12_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_12_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_12_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_12_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_12_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_12_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_12_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_entries_barrier_12_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_12_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_12_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_12_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_12_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_12_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_12_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_12_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_12_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_12_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_12_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_12_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_12_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_entries_barrier_12_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_normal_entries_barrier_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_normal_entries_barrier_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_normal_entries_barrier_1_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_1_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_1_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_1_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_1_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_1_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_1_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_1_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_1_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_1_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_1_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_1_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_1_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_1_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_normal_entries_barrier_1_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_1_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_1_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_1_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_1_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_1_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_1_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_1_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_1_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_1_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_1_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_1_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_1_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_1_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_normal_entries_barrier_2_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_2_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_2_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_2_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_2_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_2_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_2_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_2_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_2_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_2_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_2_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_2_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_2_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_2_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_normal_entries_barrier_2_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_2_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_2_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_2_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_2_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_2_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_2_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_2_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_2_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_2_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_2_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_2_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_2_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_2_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_normal_entries_barrier_3_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_3_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_3_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_3_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_3_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_3_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_3_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_3_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_3_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_3_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_3_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_3_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_3_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_3_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_normal_entries_barrier_3_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_3_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_3_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_3_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_3_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_3_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_3_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_3_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_3_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_3_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_3_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_3_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_3_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_3_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_normal_entries_barrier_4_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_4_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_4_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_4_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_4_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_4_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_4_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_4_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_4_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_4_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_4_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_4_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_4_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_4_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_normal_entries_barrier_4_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_4_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_4_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_4_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_4_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_4_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_4_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_4_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_4_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_4_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_4_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_4_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_4_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_4_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_normal_entries_barrier_5_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_5_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_5_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_5_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_5_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_5_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_5_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_5_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_5_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_5_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_5_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_5_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_5_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_5_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_normal_entries_barrier_5_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_5_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_5_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_5_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_5_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_5_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_5_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_5_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_5_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_5_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_5_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_5_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_5_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_5_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_normal_entries_barrier_6_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_6_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_6_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_6_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_6_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_6_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_6_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_6_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_6_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_6_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_6_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_6_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_6_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_6_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_normal_entries_barrier_6_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_6_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_6_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_6_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_6_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_6_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_6_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_6_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_6_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_6_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_6_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_6_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_6_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_6_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_normal_entries_barrier_7_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_7_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_7_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_7_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_7_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_7_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_7_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_7_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_7_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_7_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_7_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_7_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_7_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_7_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_normal_entries_barrier_7_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_7_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_7_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_7_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_7_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_7_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_7_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_7_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_7_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_7_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_7_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_7_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_7_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_7_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_normal_entries_barrier_8_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_8_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_8_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_8_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_8_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_8_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_8_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_8_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_8_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_8_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_8_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_8_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_8_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_8_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_normal_entries_barrier_8_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_8_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_8_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_8_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_8_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_8_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_8_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_8_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_8_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_8_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_8_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_8_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_8_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_8_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_normal_entries_barrier_9_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_9_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_9_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_9_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_9_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_9_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_9_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_9_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_9_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_9_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_9_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_9_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_9_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_9_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_normal_entries_barrier_9_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_9_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_9_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_9_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_9_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_9_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_9_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_9_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_9_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_9_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_9_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_9_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_9_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_9_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_normal_entries_barrier_10_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_10_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_10_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_10_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_10_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_10_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_10_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_10_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_10_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_10_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_10_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_10_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_10_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_10_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_normal_entries_barrier_10_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_10_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_10_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_10_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_10_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_10_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_10_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_10_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_10_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_10_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_10_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_10_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_10_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_10_io_y_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_normal_entries_barrier_11_io_x_ppn; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_11_io_x_u; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_11_io_x_ae; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_11_io_x_sw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_11_io_x_sx; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_11_io_x_sr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_11_io_x_pw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_11_io_x_px; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_11_io_x_pr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_11_io_x_ppp; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_11_io_x_pal; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_11_io_x_paa; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_11_io_x_eff; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_11_io_x_c; // @[package.scala 236:25]
  wire [19:0] pma_checker_normal_entries_barrier_11_io_y_ppn; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_11_io_y_u; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_11_io_y_ae; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_11_io_y_sw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_11_io_y_sx; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_11_io_y_sr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_11_io_y_pw; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_11_io_y_px; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_11_io_y_pr; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_11_io_y_ppp; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_11_io_y_pal; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_11_io_y_paa; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_11_io_y_eff; // @[package.scala 236:25]
  wire  pma_checker_normal_entries_barrier_11_io_y_c; // @[package.scala 236:25]
  wire  lfsr_prng_clock; // @[PRNG.scala 82:22]
  wire  lfsr_prng_reset; // @[PRNG.scala 82:22]
  wire  lfsr_prng_io_increment; // @[PRNG.scala 82:22]
  wire  lfsr_prng_io_out_0; // @[PRNG.scala 82:22]
  wire  lfsr_prng_io_out_1; // @[PRNG.scala 82:22]
  wire  lfsr_prng_io_out_2; // @[PRNG.scala 82:22]
  wire  lfsr_prng_io_out_3; // @[PRNG.scala 82:22]
  wire  lfsr_prng_io_out_4; // @[PRNG.scala 82:22]
  wire  lfsr_prng_io_out_5; // @[PRNG.scala 82:22]
  wire  lfsr_prng_io_out_6; // @[PRNG.scala 82:22]
  wire  lfsr_prng_io_out_7; // @[PRNG.scala 82:22]
  wire  lfsr_prng_io_out_8; // @[PRNG.scala 82:22]
  wire  lfsr_prng_io_out_9; // @[PRNG.scala 82:22]
  wire  lfsr_prng_io_out_10; // @[PRNG.scala 82:22]
  wire  lfsr_prng_io_out_11; // @[PRNG.scala 82:22]
  wire  lfsr_prng_io_out_12; // @[PRNG.scala 82:22]
  wire  lfsr_prng_io_out_13; // @[PRNG.scala 82:22]
  wire  lfsr_prng_io_out_14; // @[PRNG.scala 82:22]
  wire  lfsr_prng_io_out_15; // @[PRNG.scala 82:22]
  wire  metaArb_io_in_0_valid;
  wire [39:0] metaArb_io_in_0_bits_addr;
  wire [5:0] metaArb_io_in_0_bits_idx;
  wire [21:0] metaArb_io_in_0_bits_data;
  wire  metaArb_io_in_2_valid;
  wire [39:0] metaArb_io_in_2_bits_addr;
  wire [5:0] metaArb_io_in_2_bits_idx;
  wire [3:0] metaArb_io_in_2_bits_way_en;
  wire [21:0] metaArb_io_in_2_bits_data;
  wire  metaArb_io_in_3_valid;
  wire [39:0] metaArb_io_in_3_bits_addr;
  wire [5:0] metaArb_io_in_3_bits_idx;
  wire [3:0] metaArb_io_in_3_bits_way_en;
  wire [21:0] metaArb_io_in_3_bits_data;
  wire  metaArb_io_in_4_ready;
  wire  metaArb_io_in_4_valid;
  wire [39:0] metaArb_io_in_4_bits_addr;
  wire [5:0] metaArb_io_in_4_bits_idx;
  wire [3:0] metaArb_io_in_4_bits_way_en;
  wire [21:0] metaArb_io_in_4_bits_data;
  wire [39:0] metaArb_io_in_5_bits_addr;
  wire [5:0] metaArb_io_in_5_bits_idx;
  wire  metaArb_io_in_6_ready;
  wire  metaArb_io_in_6_valid;
  wire [39:0] metaArb_io_in_6_bits_addr;
  wire [5:0] metaArb_io_in_6_bits_idx;
  wire [3:0] metaArb_io_in_6_bits_way_en;
  wire [21:0] metaArb_io_in_6_bits_data;
  wire  metaArb_io_in_7_ready;
  wire  metaArb_io_in_7_valid;
  wire [39:0] metaArb_io_in_7_bits_addr;
  wire [5:0] metaArb_io_in_7_bits_idx;
  wire [3:0] metaArb_io_in_7_bits_way_en;
  wire [21:0] metaArb_io_in_7_bits_data;
  wire  metaArb_io_out_valid;
  wire  metaArb_io_out_bits_write;
  wire [39:0] metaArb_io_out_bits_addr;
  wire [5:0] metaArb_io_out_bits_idx;
  wire [3:0] metaArb_io_out_bits_way_en;
  wire [21:0] metaArb_io_out_bits_data;
  wire [21:0] metaArb__GEN_1 = metaArb_io_in_6_valid ? metaArb_io_in_6_bits_data : metaArb_io_in_7_bits_data; // @[Arbiter.scala 126:27 Arbiter.scala 128:19 Arbiter.scala 124:15]
  wire [3:0] metaArb__GEN_2 = metaArb_io_in_6_valid ? metaArb_io_in_6_bits_way_en : metaArb_io_in_7_bits_way_en; // @[Arbiter.scala 126:27 Arbiter.scala 128:19 Arbiter.scala 124:15]
  wire [5:0] metaArb__GEN_3 = metaArb_io_in_6_valid ? metaArb_io_in_6_bits_idx : metaArb_io_in_7_bits_idx; // @[Arbiter.scala 126:27 Arbiter.scala 128:19 Arbiter.scala 124:15]
  wire [39:0] metaArb__GEN_4 = metaArb_io_in_6_valid ? metaArb_io_in_6_bits_addr : metaArb_io_in_7_bits_addr; // @[Arbiter.scala 126:27 Arbiter.scala 128:19 Arbiter.scala 124:15]
  wire [21:0] metaArb__GEN_13 = metaArb_io_in_4_valid ? metaArb_io_in_4_bits_data : metaArb__GEN_1; // @[Arbiter.scala 126:27 Arbiter.scala 128:19]
  wire [3:0] metaArb__GEN_14 = metaArb_io_in_4_valid ? metaArb_io_in_4_bits_way_en : metaArb__GEN_2; // @[Arbiter.scala 126:27 Arbiter.scala 128:19]
  wire [5:0] metaArb__GEN_15 = metaArb_io_in_4_valid ? metaArb_io_in_4_bits_idx : metaArb__GEN_3; // @[Arbiter.scala 126:27 Arbiter.scala 128:19]
  wire [39:0] metaArb__GEN_16 = metaArb_io_in_4_valid ? metaArb_io_in_4_bits_addr : metaArb__GEN_4; // @[Arbiter.scala 126:27 Arbiter.scala 128:19]
  wire [21:0] metaArb__GEN_19 = metaArb_io_in_3_valid ? metaArb_io_in_3_bits_data : metaArb__GEN_13; // @[Arbiter.scala 126:27 Arbiter.scala 128:19]
  wire [3:0] metaArb__GEN_20 = metaArb_io_in_3_valid ? metaArb_io_in_3_bits_way_en : metaArb__GEN_14; // @[Arbiter.scala 126:27 Arbiter.scala 128:19]
  wire [5:0] metaArb__GEN_21 = metaArb_io_in_3_valid ? metaArb_io_in_3_bits_idx : metaArb__GEN_15; // @[Arbiter.scala 126:27 Arbiter.scala 128:19]
  wire [39:0] metaArb__GEN_22 = metaArb_io_in_3_valid ? metaArb_io_in_3_bits_addr : metaArb__GEN_16; // @[Arbiter.scala 126:27 Arbiter.scala 128:19]
  wire  metaArb__GEN_23 = metaArb_io_in_3_valid | metaArb_io_in_4_valid; // @[Arbiter.scala 126:27 Arbiter.scala 128:19]
  wire [21:0] metaArb__GEN_25 = metaArb_io_in_2_valid ? metaArb_io_in_2_bits_data : metaArb__GEN_19; // @[Arbiter.scala 126:27 Arbiter.scala 128:19]
  wire [3:0] metaArb__GEN_26 = metaArb_io_in_2_valid ? metaArb_io_in_2_bits_way_en : metaArb__GEN_20; // @[Arbiter.scala 126:27 Arbiter.scala 128:19]
  wire [5:0] metaArb__GEN_27 = metaArb_io_in_2_valid ? metaArb_io_in_2_bits_idx : metaArb__GEN_21; // @[Arbiter.scala 126:27 Arbiter.scala 128:19]
  wire [39:0] metaArb__GEN_28 = metaArb_io_in_2_valid ? metaArb_io_in_2_bits_addr : metaArb__GEN_22; // @[Arbiter.scala 126:27 Arbiter.scala 128:19]
  wire  metaArb__GEN_29 = metaArb_io_in_2_valid | metaArb__GEN_23; // @[Arbiter.scala 126:27 Arbiter.scala 128:19]
  wire  metaArb__grant_T_1 = metaArb_io_in_0_valid | metaArb_io_in_2_valid; // @[Arbiter.scala 31:68]
  wire  metaArb__grant_T_2 = metaArb__grant_T_1 | metaArb_io_in_3_valid; // @[Arbiter.scala 31:68]
  wire  metaArb__grant_T_3 = metaArb__grant_T_2 | metaArb_io_in_4_valid; // @[Arbiter.scala 31:68]
  wire  metaArb__grant_T_5 = metaArb__grant_T_3 | metaArb_io_in_6_valid; // @[Arbiter.scala 31:68]
  wire  metaArb_grant_7 = ~metaArb__grant_T_5; // @[Arbiter.scala 31:78]
  wire  metaArb__io_out_valid_T = ~metaArb_grant_7; // @[Arbiter.scala 135:19]
  wire [5:0] tag_array_RW0_addr; // @[DescribedSRAM.scala 23:26]
  wire  tag_array_RW0_en; // @[DescribedSRAM.scala 23:26]
  wire  tag_array_RW0_clk; // @[DescribedSRAM.scala 23:26]
  wire  tag_array_RW0_wmode; // @[DescribedSRAM.scala 23:26]
  wire [21:0] tag_array_RW0_wdata_0; // @[DescribedSRAM.scala 23:26]
  wire [21:0] tag_array_RW0_wdata_1; // @[DescribedSRAM.scala 23:26]
  wire [21:0] tag_array_RW0_wdata_2; // @[DescribedSRAM.scala 23:26]
  wire [21:0] tag_array_RW0_wdata_3; // @[DescribedSRAM.scala 23:26]
  wire [21:0] tag_array_RW0_rdata_0; // @[DescribedSRAM.scala 23:26]
  wire [21:0] tag_array_RW0_rdata_1; // @[DescribedSRAM.scala 23:26]
  wire [21:0] tag_array_RW0_rdata_2; // @[DescribedSRAM.scala 23:26]
  wire [21:0] tag_array_RW0_rdata_3; // @[DescribedSRAM.scala 23:26]
  wire  tag_array_RW0_wmask_0; // @[DescribedSRAM.scala 23:26]
  wire  tag_array_RW0_wmask_1; // @[DescribedSRAM.scala 23:26]
  wire  tag_array_RW0_wmask_2; // @[DescribedSRAM.scala 23:26]
  wire  tag_array_RW0_wmask_3; // @[DescribedSRAM.scala 23:26]
  wire  data_clock; // @[DCache.scala 130:20]
  wire  data_io_req_valid; // @[DCache.scala 130:20]
  wire [11:0] data_io_req_bits_addr; // @[DCache.scala 130:20]
  wire  data_io_req_bits_write; // @[DCache.scala 130:20]
  wire [63:0] data_io_req_bits_wdata; // @[DCache.scala 130:20]
  wire [7:0] data_io_req_bits_eccMask; // @[DCache.scala 130:20]
  wire [3:0] data_io_req_bits_way_en; // @[DCache.scala 130:20]
  wire [63:0] data_io_resp_0; // @[DCache.scala 130:20]
  wire [63:0] data_io_resp_1; // @[DCache.scala 130:20]
  wire [63:0] data_io_resp_2; // @[DCache.scala 130:20]
  wire [63:0] data_io_resp_3; // @[DCache.scala 130:20]
  wire  dataArb_io_in_0_valid;
  wire [11:0] dataArb_io_in_0_bits_addr;
  wire  dataArb_io_in_0_bits_write;
  wire [63:0] dataArb_io_in_0_bits_wdata;
  wire [7:0] dataArb_io_in_0_bits_eccMask;
  wire [3:0] dataArb_io_in_0_bits_way_en;
  wire  dataArb_io_in_1_ready;
  wire  dataArb_io_in_1_valid;
  wire [11:0] dataArb_io_in_1_bits_addr;
  wire  dataArb_io_in_1_bits_write;
  wire [63:0] dataArb_io_in_1_bits_wdata;
  wire [3:0] dataArb_io_in_1_bits_way_en;
  wire  dataArb_io_in_2_ready;
  wire  dataArb_io_in_2_valid;
  wire [11:0] dataArb_io_in_2_bits_addr;
  wire [63:0] dataArb_io_in_2_bits_wdata;
  wire  dataArb_io_in_3_ready;
  wire  dataArb_io_in_3_valid;
  wire [11:0] dataArb_io_in_3_bits_addr;
  wire [63:0] dataArb_io_in_3_bits_wdata;
  wire  dataArb_io_out_valid;
  wire [11:0] dataArb_io_out_bits_addr;
  wire  dataArb_io_out_bits_write;
  wire [63:0] dataArb_io_out_bits_wdata;
  wire [7:0] dataArb_io_out_bits_eccMask;
  wire [3:0] dataArb_io_out_bits_way_en;
  wire [63:0] dataArb__GEN_4 = dataArb_io_in_2_valid ? dataArb_io_in_2_bits_wdata : dataArb_io_in_3_bits_wdata; // @[Arbiter.scala 126:27 Arbiter.scala 128:19 Arbiter.scala 124:15]
  wire [11:0] dataArb__GEN_6 = dataArb_io_in_2_valid ? dataArb_io_in_2_bits_addr : dataArb_io_in_3_bits_addr; // @[Arbiter.scala 126:27 Arbiter.scala 128:19 Arbiter.scala 124:15]
  wire [3:0] dataArb__GEN_8 = dataArb_io_in_1_valid ? dataArb_io_in_1_bits_way_en : 4'hf; // @[Arbiter.scala 126:27 Arbiter.scala 128:19]
  wire [63:0] dataArb__GEN_11 = dataArb_io_in_1_valid ? dataArb_io_in_1_bits_wdata : dataArb__GEN_4; // @[Arbiter.scala 126:27 Arbiter.scala 128:19]
  wire  dataArb__GEN_12 = dataArb_io_in_1_valid & dataArb_io_in_1_bits_write; // @[Arbiter.scala 126:27 Arbiter.scala 128:19]
  wire [11:0] dataArb__GEN_13 = dataArb_io_in_1_valid ? dataArb_io_in_1_bits_addr : dataArb__GEN_6; // @[Arbiter.scala 126:27 Arbiter.scala 128:19]
  wire  dataArb__grant_T = dataArb_io_in_0_valid | dataArb_io_in_1_valid; // @[Arbiter.scala 31:68]
  wire  dataArb__grant_T_1 = dataArb__grant_T | dataArb_io_in_2_valid; // @[Arbiter.scala 31:68]
  wire  dataArb_grant_3 = ~dataArb__grant_T_1; // @[Arbiter.scala 31:78]
  wire  dataArb__io_out_valid_T = ~dataArb_grant_3; // @[Arbiter.scala 135:19]
  wire [7:0] amoalu_io_mask; // @[DCache.scala 881:26]
  wire [4:0] amoalu_io_cmd; // @[DCache.scala 881:26]
  wire [63:0] amoalu_io_lhs; // @[DCache.scala 881:26]
  wire [63:0] amoalu_io_rhs; // @[DCache.scala 881:26]
  wire [63:0] amoalu_io_out; // @[DCache.scala 881:26]
  wire [7:0] lfsr_left = {lfsr_prng_io_out_7,lfsr_prng_io_out_6,lfsr_prng_io_out_5,lfsr_prng_io_out_4,lfsr_prng_io_out_3
    ,lfsr_prng_io_out_2,lfsr_prng_io_out_1,lfsr_prng_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] lfsr = {lfsr_prng_io_out_15,lfsr_prng_io_out_14,lfsr_prng_io_out_13,lfsr_prng_io_out_12,
    lfsr_prng_io_out_11,lfsr_prng_io_out_10,lfsr_prng_io_out_9,lfsr_prng_io_out_8,lfsr_left}; // @[PRNG.scala 86:17]
  wire  s1_valid_x9 = io_cpu_req_ready & io_cpu_req_valid; // @[Decoupled.scala 40:37]
  reg  s1_valid; // @[DCache.scala 159:21]
  reg [2:0] blockProbeAfterGrantCount; // @[DCache.scala 611:38]
  wire  _block_probe_for_core_progress_T = blockProbeAfterGrantCount > 3'h0; // @[DCache.scala 709:65]
  reg [6:0] lrscCount; // @[DCache.scala 423:22]
  wire  lrscValid = lrscCount > 7'h3; // @[DCache.scala 424:29]
  wire  block_probe_for_core_progress = (blockProbeAfterGrantCount > 3'h0) | lrscValid; // @[DCache.scala 709:69]
  reg  s1_probe; // @[DCache.scala 160:21]
  reg  s2_probe; // @[DCache.scala 285:21]
  reg [2:0] release_state; // @[DCache.scala 199:26]
  wire  releaseInFlight = (s1_probe | s2_probe) | (release_state != 3'h0); // @[DCache.scala 286:46]
  reg  release_ack_wait; // @[DCache.scala 197:29]
  reg [31:0] release_ack_addr; // @[DCache.scala 198:29]
  wire [31:0] _block_probe_for_pending_release_ack_T = auto_out_b_bits_address ^ release_ack_addr; // @[DCache.scala 710:88]
  wire  block_probe_for_pending_release_ack = release_ack_wait & ((_block_probe_for_pending_release_ack_T[11:6]) == 6'h0
    ); // @[DCache.scala 710:62]
  reg  grantInProgress; // @[DCache.scala 610:28]
  wire  block_probe_for_ordering = (releaseInFlight | block_probe_for_pending_release_ack) | grantInProgress; // @[DCache.scala 711:89]
  reg  s2_valid; // @[DCache.scala 283:21]
  wire  tl_out__b_ready = metaArb_io_in_6_ready & (~(((block_probe_for_core_progress | block_probe_for_ordering) |
    s1_valid) | s2_valid)); // @[DCache.scala 713:44]
  wire  s1_probe_x12 = tl_out__b_ready & auto_out_b_valid; // @[Decoupled.scala 40:37]
  reg [1:0] probe_bits_param; // @[Reg.scala 15:16]
  reg [3:0] probe_bits_size; // @[Reg.scala 15:16]
  reg  probe_bits_source; // @[Reg.scala 15:16]
  reg [31:0] probe_bits_address; // @[Reg.scala 15:16]
  wire  s1_valid_masked = s1_valid & (~io_cpu_s1_kill); // @[DCache.scala 163:34]
  reg [1:0] s2_probe_state_state; // @[Reg.scala 15:16]
  wire [3:0] _T_83 = {probe_bits_param,s2_probe_state_state}; // @[Cat.scala 29:58]
  wire  _T_140 = 4'h3 == _T_83; // @[Misc.scala 55:20]
  wire  _T_136 = 4'h2 == _T_83; // @[Misc.scala 55:20]
  wire  _T_132 = 4'h1 == _T_83; // @[Misc.scala 55:20]
  wire  _T_128 = 4'h0 == _T_83; // @[Misc.scala 55:20]
  wire  _T_124 = 4'h7 == _T_83; // @[Misc.scala 55:20]
  wire  _T_120 = 4'h6 == _T_83; // @[Misc.scala 55:20]
  wire  _T_116 = 4'h5 == _T_83; // @[Misc.scala 55:20]
  wire  _T_112 = 4'h4 == _T_83; // @[Misc.scala 55:20]
  wire  _T_108 = 4'hb == _T_83; // @[Misc.scala 55:20]
  wire  _T_104 = 4'ha == _T_83; // @[Misc.scala 55:20]
  wire  _T_100 = 4'h9 == _T_83; // @[Misc.scala 55:20]
  wire  _T_96 = 4'h8 == _T_83; // @[Misc.scala 55:20]
  wire  _T_113 = _T_112 ? 1'h0 : _T_108; // @[Misc.scala 37:9]
  wire  _T_117 = _T_116 ? 1'h0 : _T_113; // @[Misc.scala 37:9]
  wire  _T_121 = _T_120 ? 1'h0 : _T_117; // @[Misc.scala 37:9]
  wire  _T_129 = _T_128 ? 1'h0 : _T_124 | _T_121; // @[Misc.scala 37:9]
  wire  _T_133 = _T_132 ? 1'h0 : _T_129; // @[Misc.scala 37:9]
  wire  _T_137 = _T_136 ? 1'h0 : _T_133; // @[Misc.scala 37:9]
  wire  s2_prb_ack_data = _T_140 | _T_137; // @[Misc.scala 37:9]
  wire  _T_268 = s2_probe_state_state > 2'h0; // @[Metadata.scala 50:45]
  reg [8:0] counter_1; // @[Edges.scala 230:27]
  wire  _T_273 = release_state == 3'h1; // @[package.scala 15:47]
  wire  _T_274 = release_state == 3'h6; // @[package.scala 15:47]
  wire  _T_275 = _T_273 | _T_274; // @[package.scala 64:59]
  wire  _T_272 = release_state == 3'h2; // @[DCache.scala 779:25]
  wire  _T_271 = release_state == 3'h3; // @[DCache.scala 774:25]
  wire [2:0] _GEN_314 = _T_272 ? 3'h5 : 3'h4; // @[DCache.scala 779:48 DCache.scala 780:21]
  wire [2:0] tl_out__c_bits_opcode = _T_275 ? 3'h7 : _GEN_314; // @[DCache.scala 783:81 DCache.scala 784:21]
  wire  beats1_opdata_1 = tl_out__c_bits_opcode[0]; // @[Edges.scala 103:36]
  wire [3:0] tl_out__c_bits_size = _T_275 ? 4'h6 : probe_bits_size; // @[DCache.scala 783:81 DCache.scala 784:21]
  wire [26:0] _beats1_decode_T_5 = 27'hfff << tl_out__c_bits_size; // @[package.scala 212:77]
  wire [11:0] _beats1_decode_T_7 = ~(_beats1_decode_T_5[11:0]); // @[package.scala 212:46]
  wire [8:0] beats1_decode_1 = _beats1_decode_T_7[11:3]; // @[Edges.scala 221:59]
  wire [8:0] beats1_1 = beats1_opdata_1 ? beats1_decode_1 : 9'h0; // @[Edges.scala 222:14]
  wire  c_last = (counter_1 == 9'h1) | (beats1_1 == 9'h0); // @[Edges.scala 233:37]
  wire  _T_270 = release_state == 3'h5; // @[DCache.scala 770:25]
  reg  s2_release_data_valid; // @[DCache.scala 724:34]
  wire  c_first = counter_1 == 9'h0; // @[Edges.scala 232:25]
  wire  _tl_out_c_valid_T_2 = s2_release_data_valid & (~(c_first & release_ack_wait)); // @[DCache.scala 732:43]
  wire  _GEN_263 = s2_prb_ack_data ? _tl_out_c_valid_T_2 : 1'h1; // @[DCache.scala 748:36 DCache.scala 732:18]
  wire  _GEN_284 = s2_probe ? _GEN_263 : _tl_out_c_valid_T_2; // @[DCache.scala 744:21 DCache.scala 732:18]
  wire  _GEN_301 = _T_270 | _GEN_284; // @[DCache.scala 770:47 DCache.scala 771:22]
  wire  tl_out__c_valid = _T_271 | _GEN_301; // @[DCache.scala 774:48 DCache.scala 775:22]
  wire  _T_262 = auto_out_c_ready & tl_out__c_valid; // @[Decoupled.scala 40:37]
  wire  releaseDone = c_last & _T_262; // @[Edges.scala 234:22]
  wire  _probeNack_T = ~releaseDone; // @[DCache.scala 756:22]
  wire  _GEN_261 = _T_268 | _probeNack_T; // @[DCache.scala 750:45 DCache.scala 756:19]
  wire  probeNack = s2_prb_ack_data | _GEN_261; // @[DCache.scala 748:36]
  reg [4:0] s1_req_cmd; // @[Reg.scala 15:16]
  wire  _s1_read_T_3 = s1_req_cmd == 5'h7; // @[Consts.scala 82:65]
  wire  _s1_read_T_5 = s1_req_cmd == 5'h4; // @[package.scala 15:47]
  wire  _s1_read_T_6 = s1_req_cmd == 5'h9; // @[package.scala 15:47]
  wire  _s1_read_T_7 = s1_req_cmd == 5'ha; // @[package.scala 15:47]
  wire  _s1_read_T_8 = s1_req_cmd == 5'hb; // @[package.scala 15:47]
  wire  _s1_read_T_11 = ((_s1_read_T_5 | _s1_read_T_6) | _s1_read_T_7) | _s1_read_T_8; // @[package.scala 64:59]
  wire  _s1_read_T_12 = s1_req_cmd == 5'h8; // @[package.scala 15:47]
  wire  _s1_read_T_13 = s1_req_cmd == 5'hc; // @[package.scala 15:47]
  wire  _s1_read_T_14 = s1_req_cmd == 5'hd; // @[package.scala 15:47]
  wire  _s1_read_T_15 = s1_req_cmd == 5'he; // @[package.scala 15:47]
  wire  _s1_read_T_16 = s1_req_cmd == 5'hf; // @[package.scala 15:47]
  wire  _s1_read_T_20 = (((_s1_read_T_12 | _s1_read_T_13) | _s1_read_T_14) | _s1_read_T_15) | _s1_read_T_16; // @[package.scala 64:59]
  wire  _s1_read_T_21 = _s1_read_T_11 | _s1_read_T_20; // @[Consts.scala 80:44]
  wire  s1_read = (((s1_req_cmd == 5'h0) | (s1_req_cmd == 5'h6)) | (s1_req_cmd == 5'h7)) | _s1_read_T_21; // @[Consts.scala 82:75]
  reg [4:0] s2_req_cmd; // @[DCache.scala 291:19]
  wire  _s2_write_T_1 = s2_req_cmd == 5'h11; // @[Consts.scala 83:49]
  wire  _s2_write_T_3 = s2_req_cmd == 5'h7; // @[Consts.scala 83:66]
  wire  _s2_write_T_5 = s2_req_cmd == 5'h4; // @[package.scala 15:47]
  wire  _s2_write_T_6 = s2_req_cmd == 5'h9; // @[package.scala 15:47]
  wire  _s2_write_T_7 = s2_req_cmd == 5'ha; // @[package.scala 15:47]
  wire  _s2_write_T_8 = s2_req_cmd == 5'hb; // @[package.scala 15:47]
  wire  _s2_write_T_11 = ((_s2_write_T_5 | _s2_write_T_6) | _s2_write_T_7) | _s2_write_T_8; // @[package.scala 64:59]
  wire  _s2_write_T_12 = s2_req_cmd == 5'h8; // @[package.scala 15:47]
  wire  _s2_write_T_13 = s2_req_cmd == 5'hc; // @[package.scala 15:47]
  wire  _s2_write_T_14 = s2_req_cmd == 5'hd; // @[package.scala 15:47]
  wire  _s2_write_T_15 = s2_req_cmd == 5'he; // @[package.scala 15:47]
  wire  _s2_write_T_16 = s2_req_cmd == 5'hf; // @[package.scala 15:47]
  wire  _s2_write_T_20 = (((_s2_write_T_12 | _s2_write_T_13) | _s2_write_T_14) | _s2_write_T_15) | _s2_write_T_16; // @[package.scala 64:59]
  wire  _s2_write_T_21 = _s2_write_T_11 | _s2_write_T_20; // @[Consts.scala 80:44]
  wire  s2_write = (((s2_req_cmd == 5'h1) | (s2_req_cmd == 5'h11)) | (s2_req_cmd == 5'h7)) | _s2_write_T_21; // @[Consts.scala 83:76]
  reg  pstore1_held; // @[DCache.scala 455:25]
  wire  pstore1_valid_likely = (s2_valid & s2_write) | pstore1_held; // @[DCache.scala 456:51]
  reg [39:0] pstore1_addr; // @[Reg.scala 15:16]
  reg [39:0] s1_req_addr; // @[Reg.scala 15:16]
  wire  _s1_write_T_1 = s1_req_cmd == 5'h11; // @[Consts.scala 83:49]
  wire  s1_write = (((s1_req_cmd == 5'h1) | (s1_req_cmd == 5'h11)) | _s1_read_T_3) | _s1_read_T_21; // @[Consts.scala 83:76]
  reg [7:0] pstore1_mask; // @[Reg.scala 15:16]
  wire  s1_hazard_right_right_right = |(pstore1_mask[7]); // @[DCache.scala 1076:66]
  wire  s1_hazard_right_right_left = |(pstore1_mask[6]); // @[DCache.scala 1076:66]
  wire  s1_hazard_right_left_right = |(pstore1_mask[5]); // @[DCache.scala 1076:66]
  wire  s1_hazard_right_left_left = |(pstore1_mask[4]); // @[DCache.scala 1076:66]
  wire  s1_hazard_left_right_right = |(pstore1_mask[3]); // @[DCache.scala 1076:66]
  wire  s1_hazard_left_right_left = |(pstore1_mask[2]); // @[DCache.scala 1076:66]
  wire  s1_hazard_left_left_right = |(pstore1_mask[1]); // @[DCache.scala 1076:66]
  wire  s1_hazard_left_left_left = |(pstore1_mask[0]); // @[DCache.scala 1076:66]
  wire [7:0] _s1_hazard_T_11 = {s1_hazard_right_right_right,s1_hazard_right_right_left,s1_hazard_right_left_right,
    s1_hazard_right_left_left,s1_hazard_left_right_right,s1_hazard_left_right_left,s1_hazard_left_left_right,
    s1_hazard_left_left_left}; // @[Cat.scala 29:58]
  wire  s1_hazard_right_right_right_1 = _s1_hazard_T_11[7]; // @[Bitwise.scala 26:51]
  wire  s1_hazard_right_right_left_1 = _s1_hazard_T_11[6]; // @[Bitwise.scala 26:51]
  wire  s1_hazard_right_left_right_1 = _s1_hazard_T_11[5]; // @[Bitwise.scala 26:51]
  wire  s1_hazard_right_left_left_1 = _s1_hazard_T_11[4]; // @[Bitwise.scala 26:51]
  wire  s1_hazard_left_right_right_1 = _s1_hazard_T_11[3]; // @[Bitwise.scala 26:51]
  wire  s1_hazard_left_right_left_1 = _s1_hazard_T_11[2]; // @[Bitwise.scala 26:51]
  wire  s1_hazard_left_left_right_1 = _s1_hazard_T_11[1]; // @[Bitwise.scala 26:51]
  wire  s1_hazard_left_left_left_1 = _s1_hazard_T_11[0]; // @[Bitwise.scala 26:51]
  wire [7:0] _s1_hazard_T_12 = {s1_hazard_right_right_right_1,s1_hazard_right_right_left_1,s1_hazard_right_left_right_1,
    s1_hazard_right_left_left_1,s1_hazard_left_right_right_1,s1_hazard_left_right_left_1,s1_hazard_left_left_right_1,
    s1_hazard_left_left_left_1}; // @[Cat.scala 29:58]
  reg [1:0] s1_req_size; // @[Reg.scala 15:16]
  wire  s1_mask_xwr_right = (s1_req_addr[0]) | (s1_req_size >= 2'h1); // @[AMOALU.scala 17:46]
  wire  s1_mask_xwr_left = s1_req_addr[0] ? 1'h0 : 1'h1; // @[AMOALU.scala 18:22]
  wire [1:0] _s1_mask_xwr_T = {s1_mask_xwr_right,s1_mask_xwr_left}; // @[Cat.scala 29:58]
  wire [1:0] _s1_mask_xwr_upper_T_5 = s1_req_addr[1] ? _s1_mask_xwr_T : 2'h0; // @[AMOALU.scala 17:22]
  wire [1:0] _s1_mask_xwr_upper_T_7 = s1_req_size >= 2'h2 ? 2'h3 : 2'h0; // @[AMOALU.scala 17:51]
  wire [1:0] s1_mask_xwr_right_1 = _s1_mask_xwr_upper_T_5 | _s1_mask_xwr_upper_T_7; // @[AMOALU.scala 17:46]
  wire [1:0] s1_mask_xwr_left_1 = s1_req_addr[1] ? 2'h0 : _s1_mask_xwr_T; // @[AMOALU.scala 18:22]
  wire [3:0] _s1_mask_xwr_T_1 = {s1_mask_xwr_right_1,s1_mask_xwr_left_1}; // @[Cat.scala 29:58]
  wire [3:0] _s1_mask_xwr_upper_T_9 = s1_req_addr[2] ? _s1_mask_xwr_T_1 : 4'h0; // @[AMOALU.scala 17:22]
  wire [3:0] _s1_mask_xwr_upper_T_11 = s1_req_size >= 2'h3 ? 4'hf : 4'h0; // @[AMOALU.scala 17:51]
  wire [3:0] s1_mask_xwr_right_2 = _s1_mask_xwr_upper_T_9 | _s1_mask_xwr_upper_T_11; // @[AMOALU.scala 17:46]
  wire [3:0] s1_mask_xwr_left_2 = s1_req_addr[2] ? 4'h0 : _s1_mask_xwr_T_1; // @[AMOALU.scala 18:22]
  wire [7:0] s1_mask_xwr = {s1_mask_xwr_right_2,s1_mask_xwr_left_2}; // @[Cat.scala 29:58]
  wire  s1_hazard_right_right_right_2 = |(s1_mask_xwr[7]); // @[DCache.scala 1076:66]
  wire  s1_hazard_right_right_left_2 = |(s1_mask_xwr[6]); // @[DCache.scala 1076:66]
  wire  s1_hazard_right_left_right_2 = |(s1_mask_xwr[5]); // @[DCache.scala 1076:66]
  wire  s1_hazard_right_left_left_2 = |(s1_mask_xwr[4]); // @[DCache.scala 1076:66]
  wire  s1_hazard_left_right_right_2 = |(s1_mask_xwr[3]); // @[DCache.scala 1076:66]
  wire  s1_hazard_left_right_left_2 = |(s1_mask_xwr[2]); // @[DCache.scala 1076:66]
  wire  s1_hazard_left_left_right_2 = |(s1_mask_xwr[1]); // @[DCache.scala 1076:66]
  wire  s1_hazard_left_left_left_2 = |(s1_mask_xwr[0]); // @[DCache.scala 1076:66]
  wire [7:0] _s1_hazard_T_21 = {s1_hazard_right_right_right_2,s1_hazard_right_right_left_2,s1_hazard_right_left_right_2,
    s1_hazard_right_left_left_2,s1_hazard_left_right_right_2,s1_hazard_left_right_left_2,s1_hazard_left_left_right_2,
    s1_hazard_left_left_left_2}; // @[Cat.scala 29:58]
  wire  s1_hazard_right_right_right_3 = _s1_hazard_T_21[7]; // @[Bitwise.scala 26:51]
  wire  s1_hazard_right_right_left_3 = _s1_hazard_T_21[6]; // @[Bitwise.scala 26:51]
  wire  s1_hazard_right_left_right_3 = _s1_hazard_T_21[5]; // @[Bitwise.scala 26:51]
  wire  s1_hazard_right_left_left_3 = _s1_hazard_T_21[4]; // @[Bitwise.scala 26:51]
  wire  s1_hazard_left_right_right_3 = _s1_hazard_T_21[3]; // @[Bitwise.scala 26:51]
  wire  s1_hazard_left_right_left_3 = _s1_hazard_T_21[2]; // @[Bitwise.scala 26:51]
  wire  s1_hazard_left_left_right_3 = _s1_hazard_T_21[1]; // @[Bitwise.scala 26:51]
  wire  s1_hazard_left_left_left_3 = _s1_hazard_T_21[0]; // @[Bitwise.scala 26:51]
  wire [7:0] _s1_hazard_T_22 = {s1_hazard_right_right_right_3,s1_hazard_right_right_left_3,s1_hazard_right_left_right_3,
    s1_hazard_right_left_left_3,s1_hazard_left_right_right_3,s1_hazard_left_right_left_3,s1_hazard_left_left_right_3,
    s1_hazard_left_left_left_3}; // @[Cat.scala 29:58]
  wire [7:0] _s1_hazard_T_23 = _s1_hazard_T_12 & _s1_hazard_T_22; // @[DCache.scala 509:38]
  wire [7:0] _s1_hazard_T_25 = pstore1_mask & s1_mask_xwr; // @[DCache.scala 509:77]
  wire  _s1_hazard_T_27 = s1_write ? |_s1_hazard_T_23 : |_s1_hazard_T_25; // @[DCache.scala 509:8]
  wire  _s1_hazard_T_28 = ((pstore1_addr[11:3]) == (s1_req_addr[11:3])) & _s1_hazard_T_27; // @[DCache.scala 508:68]
  reg  pstore2_valid; // @[DCache.scala 452:26]
  reg [39:0] pstore2_addr; // @[Reg.scala 15:16]
  reg [7:0] mask; // @[DCache.scala 482:19]
  wire  s1_hazard_right_right_right_4 = |(mask[7]); // @[DCache.scala 1076:66]
  wire  s1_hazard_right_right_left_4 = |(mask[6]); // @[DCache.scala 1076:66]
  wire  s1_hazard_right_left_right_4 = |(mask[5]); // @[DCache.scala 1076:66]
  wire  s1_hazard_right_left_left_4 = |(mask[4]); // @[DCache.scala 1076:66]
  wire  s1_hazard_left_right_right_4 = |(mask[3]); // @[DCache.scala 1076:66]
  wire  s1_hazard_left_right_left_4 = |(mask[2]); // @[DCache.scala 1076:66]
  wire  s1_hazard_left_left_right_4 = |(mask[1]); // @[DCache.scala 1076:66]
  wire  s1_hazard_left_left_left_4 = |(mask[0]); // @[DCache.scala 1076:66]
  wire [7:0] _s1_hazard_T_41 = {s1_hazard_right_right_right_4,s1_hazard_right_right_left_4,s1_hazard_right_left_right_4,
    s1_hazard_right_left_left_4,s1_hazard_left_right_right_4,s1_hazard_left_right_left_4,s1_hazard_left_left_right_4,
    s1_hazard_left_left_left_4}; // @[Cat.scala 29:58]
  wire  s1_hazard_right_right_right_5 = _s1_hazard_T_41[7]; // @[Bitwise.scala 26:51]
  wire  s1_hazard_right_right_left_5 = _s1_hazard_T_41[6]; // @[Bitwise.scala 26:51]
  wire  s1_hazard_right_left_right_5 = _s1_hazard_T_41[5]; // @[Bitwise.scala 26:51]
  wire  s1_hazard_right_left_left_5 = _s1_hazard_T_41[4]; // @[Bitwise.scala 26:51]
  wire  s1_hazard_left_right_right_5 = _s1_hazard_T_41[3]; // @[Bitwise.scala 26:51]
  wire  s1_hazard_left_right_left_5 = _s1_hazard_T_41[2]; // @[Bitwise.scala 26:51]
  wire  s1_hazard_left_left_right_5 = _s1_hazard_T_41[1]; // @[Bitwise.scala 26:51]
  wire  s1_hazard_left_left_left_5 = _s1_hazard_T_41[0]; // @[Bitwise.scala 26:51]
  wire [7:0] _s1_hazard_T_42 = {s1_hazard_right_right_right_5,s1_hazard_right_right_left_5,s1_hazard_right_left_right_5,
    s1_hazard_right_left_left_5,s1_hazard_left_right_right_5,s1_hazard_left_right_left_5,s1_hazard_left_left_right_5,
    s1_hazard_left_left_left_5}; // @[Cat.scala 29:58]
  wire [7:0] _s1_hazard_T_53 = _s1_hazard_T_42 & _s1_hazard_T_22; // @[DCache.scala 509:38]
  wire [7:0] _s1_hazard_T_55 = mask & s1_mask_xwr; // @[DCache.scala 509:77]
  wire  _s1_hazard_T_57 = s1_write ? |_s1_hazard_T_53 : |_s1_hazard_T_55; // @[DCache.scala 509:8]
  wire  _s1_hazard_T_58 = ((pstore2_addr[11:3]) == (s1_req_addr[11:3])) & _s1_hazard_T_57; // @[DCache.scala 508:68]
  wire  _s1_hazard_T_59 = pstore2_valid & _s1_hazard_T_58; // @[DCache.scala 512:21]
  wire  s1_hazard = (pstore1_valid_likely & _s1_hazard_T_28) | _s1_hazard_T_59; // @[DCache.scala 511:69]
  wire  s1_raw_hazard = s1_read & s1_hazard; // @[DCache.scala 513:31]
  wire  _T_227 = s1_valid & s1_raw_hazard; // @[DCache.scala 518:18]
  wire [5:0] _s2_valid_no_xcpt_T = {io_cpu_s2_xcpt_ma_ld,io_cpu_s2_xcpt_ma_st,io_cpu_s2_xcpt_pf_ld,io_cpu_s2_xcpt_pf_st,
    io_cpu_s2_xcpt_ae_ld,io_cpu_s2_xcpt_ae_st}; // @[DCache.scala 284:54]
  wire  s2_valid_no_xcpt = s2_valid & (~(|_s2_valid_no_xcpt_T)); // @[DCache.scala 284:35]
  reg  s2_not_nacked_in_s1; // @[DCache.scala 287:36]
  wire  s2_valid_masked = s2_valid_no_xcpt & s2_not_nacked_in_s1; // @[DCache.scala 289:42]
  wire  _c_cat_T_47 = s2_req_cmd == 5'h6; // @[Consts.scala 84:71]
  wire  c_cat_left = (s2_write | (s2_req_cmd == 5'h3)) | (s2_req_cmd == 5'h6); // @[Consts.scala 84:64]
  reg [1:0] s2_hit_state_state; // @[Reg.scala 15:16]
  wire [3:0] _T_36 = {s2_write,c_cat_left,s2_hit_state_state}; // @[Cat.scala 29:58]
  wire  _T_82 = 4'h3 == _T_36; // @[Misc.scala 48:20]
  wire  _T_79 = 4'h2 == _T_36; // @[Misc.scala 48:20]
  wire  _T_76 = 4'h1 == _T_36; // @[Misc.scala 48:20]
  wire  _T_73 = 4'h7 == _T_36; // @[Misc.scala 48:20]
  wire  _T_70 = 4'h6 == _T_36; // @[Misc.scala 48:20]
  wire  _T_67 = 4'hf == _T_36; // @[Misc.scala 48:20]
  wire  _T_64 = 4'he == _T_36; // @[Misc.scala 48:20]
  wire  _T_61 = 4'h0 == _T_36; // @[Misc.scala 48:20]
  wire  _T_58 = 4'h5 == _T_36; // @[Misc.scala 48:20]
  wire  _T_55 = 4'h4 == _T_36; // @[Misc.scala 48:20]
  wire  _T_52 = 4'hd == _T_36; // @[Misc.scala 48:20]
  wire  _T_49 = 4'hc == _T_36; // @[Misc.scala 48:20]
  wire  s2_hit = _T_82 | (_T_79 | (_T_76 | (_T_73 | (_T_70 | (_T_67 | _T_64))))); // @[Misc.scala 34:9]
  wire  s2_valid_hit_maybe_flush_pre_data_ecc_and_waw = s2_valid_masked & s2_hit; // @[DCache.scala 349:89]
  wire  s2_read = (((s2_req_cmd == 5'h0) | _c_cat_T_47) | _s2_write_T_3) | _s2_write_T_21; // @[Consts.scala 82:75]
  wire  s2_readwrite = s2_read | s2_write; // @[DCache.scala 306:30]
  wire  s2_valid_hit_pre_data_ecc_and_waw = s2_valid_hit_maybe_flush_pre_data_ecc_and_waw & s2_readwrite; // @[DCache.scala 370:89]
  wire [1:0] _T_51 = _T_49 ? 2'h1 : 2'h0; // @[Misc.scala 34:36]
  wire [1:0] _T_54 = _T_52 ? 2'h2 : _T_51; // @[Misc.scala 34:36]
  wire [1:0] _T_57 = _T_55 ? 2'h1 : _T_54; // @[Misc.scala 34:36]
  wire [1:0] _T_60 = _T_58 ? 2'h2 : _T_57; // @[Misc.scala 34:36]
  wire [1:0] _T_63 = _T_61 ? 2'h0 : _T_60; // @[Misc.scala 34:36]
  wire [1:0] _T_66 = _T_64 ? 2'h3 : _T_63; // @[Misc.scala 34:36]
  wire [1:0] _T_69 = _T_67 ? 2'h3 : _T_66; // @[Misc.scala 34:36]
  wire [1:0] _T_72 = _T_70 ? 2'h2 : _T_69; // @[Misc.scala 34:36]
  wire [1:0] _T_75 = _T_73 ? 2'h3 : _T_72; // @[Misc.scala 34:36]
  wire [1:0] _T_78 = _T_76 ? 2'h1 : _T_75; // @[Misc.scala 34:36]
  wire [1:0] _T_81 = _T_79 ? 2'h2 : _T_78; // @[Misc.scala 34:36]
  wire [1:0] s2_grow_param = _T_82 ? 2'h3 : _T_81; // @[Misc.scala 34:36]
  wire  _s2_update_meta_T = s2_hit_state_state == s2_grow_param; // @[Metadata.scala 46:46]
  wire  s2_update_meta = ~_s2_update_meta_T; // @[Metadata.scala 47:40]
  wire  _T_207 = io_cpu_s2_nack | (s2_valid_hit_pre_data_ecc_and_waw & s2_update_meta); // @[DCache.scala 397:24]
  wire  s1_readwrite = s1_read | s1_write; // @[DCache.scala 185:30]
  wire  s1_flush_line = (s1_req_cmd == 5'h5) & (s1_req_size[0]); // @[DCache.scala 187:50]
  wire  s1_cmd_uses_tlb = (s1_readwrite | s1_flush_line) | (s1_req_cmd == 5'h17); // @[DCache.scala 229:55]
  wire  _T_14 = (s1_valid & s1_cmd_uses_tlb) & tlb_io_resp_miss; // @[DCache.scala 235:58]
  wire  _GEN_118 = _T_207 | _T_14; // @[DCache.scala 397:82 DCache.scala 397:92]
  wire  _GEN_142 = _T_227 | _GEN_118; // @[DCache.scala 518:36 DCache.scala 518:46]
  wire  _GEN_282 = probeNack | _GEN_142; // @[DCache.scala 759:24 DCache.scala 759:34]
  wire  s1_nack = s2_probe ? _GEN_282 : _GEN_142; // @[DCache.scala 744:21]
  wire  _s1_valid_not_nacked_T = ~s1_nack; // @[DCache.scala 164:41]
  wire  s1_valid_not_nacked = s1_valid & (~s1_nack); // @[DCache.scala 164:38]
  wire  s0_clk_en = metaArb_io_out_valid & (~metaArb_io_out_bits_write); // @[DCache.scala 167:40]
  wire [33:0] s0_req_addr_right = metaArb_io_out_bits_addr[39:6]; // @[DCache.scala 170:47]
  wire [5:0] s0_req_addr_left = io_cpu_req_bits_addr[5:0]; // @[DCache.scala 170:84]
  wire [39:0] s0_req_addr = {s0_req_addr_right,s0_req_addr_left}; // @[Cat.scala 29:58]
  wire  _T = ~metaArb_io_in_7_ready; // @[DCache.scala 171:9]
  wire  s0_req_phys = _T | io_cpu_req_bits_phys; // @[DCache.scala 171:34 DCache.scala 171:48]
  reg [6:0] s1_req_tag; // @[Reg.scala 15:16]
  reg  s1_req_signed; // @[Reg.scala 15:16]
  reg [1:0] s1_req_dprv; // @[Reg.scala 15:16]
  reg [39:0] s1_tlb_req_vaddr; // @[Reg.scala 15:16]
  reg  s1_tlb_req_passthrough; // @[Reg.scala 15:16]
  reg [1:0] s1_tlb_req_size; // @[Reg.scala 15:16]
  reg [4:0] s1_tlb_req_cmd; // @[Reg.scala 15:16]
  wire  s1_sfence = s1_req_cmd == 5'h14; // @[DCache.scala 186:30]
  reg  cached_grant_wait; // @[DCache.scala 196:30]
  wire  inWriteback = _T_273 | _T_272; // @[package.scala 64:59]
  wire  _io_cpu_req_ready_T_1 = ~cached_grant_wait; // @[DCache.scala 203:54]
  wire  _io_cpu_req_ready_T_4 = ((release_state == 3'h0) & (~cached_grant_wait)) & _s1_valid_not_nacked_T; // @[DCache.scala 203:73]
  reg  uncachedInFlight_0; // @[DCache.scala 206:33]
  reg [39:0] uncachedReqs_0_addr; // @[DCache.scala 207:25]
  reg [6:0] uncachedReqs_0_tag; // @[DCache.scala 207:25]
  reg [1:0] uncachedReqs_0_size; // @[DCache.scala 207:25]
  reg  uncachedReqs_0_signed; // @[DCache.scala 207:25]
  wire  _s0_read_T_3 = io_cpu_req_bits_cmd == 5'h7; // @[Consts.scala 82:65]
  wire  _s0_read_T_5 = io_cpu_req_bits_cmd == 5'h4; // @[package.scala 15:47]
  wire  _s0_read_T_6 = io_cpu_req_bits_cmd == 5'h9; // @[package.scala 15:47]
  wire  _s0_read_T_7 = io_cpu_req_bits_cmd == 5'ha; // @[package.scala 15:47]
  wire  _s0_read_T_8 = io_cpu_req_bits_cmd == 5'hb; // @[package.scala 15:47]
  wire  _s0_read_T_11 = ((_s0_read_T_5 | _s0_read_T_6) | _s0_read_T_7) | _s0_read_T_8; // @[package.scala 64:59]
  wire  _s0_read_T_12 = io_cpu_req_bits_cmd == 5'h8; // @[package.scala 15:47]
  wire  _s0_read_T_13 = io_cpu_req_bits_cmd == 5'hc; // @[package.scala 15:47]
  wire  _s0_read_T_14 = io_cpu_req_bits_cmd == 5'hd; // @[package.scala 15:47]
  wire  _s0_read_T_15 = io_cpu_req_bits_cmd == 5'he; // @[package.scala 15:47]
  wire  _s0_read_T_16 = io_cpu_req_bits_cmd == 5'hf; // @[package.scala 15:47]
  wire  _s0_read_T_20 = (((_s0_read_T_12 | _s0_read_T_13) | _s0_read_T_14) | _s0_read_T_15) | _s0_read_T_16; // @[package.scala 64:59]
  wire  _s0_read_T_21 = _s0_read_T_11 | _s0_read_T_20; // @[Consts.scala 80:44]
  wire  s0_read = (((io_cpu_req_bits_cmd == 5'h0) | (io_cpu_req_bits_cmd == 5'h6)) | (io_cpu_req_bits_cmd == 5'h7)) |
    _s0_read_T_21; // @[Consts.scala 82:75]
  wire  _dataArb_io_in_3_valid_res_T = io_cpu_req_bits_cmd == 5'h1; // @[package.scala 15:47]
  wire  _dataArb_io_in_3_valid_res_T_1 = io_cpu_req_bits_cmd == 5'h3; // @[package.scala 15:47]
  wire  _dataArb_io_in_3_valid_res_T_2 = _dataArb_io_in_3_valid_res_T | _dataArb_io_in_3_valid_res_T_1; // @[package.scala 64:59]
  wire  res = ~_dataArb_io_in_3_valid_res_T_2; // @[DCache.scala 1080:15]
  wire  _dataArb_io_in_3_valid_T_24 = io_cpu_req_bits_cmd == 5'h11; // @[Consts.scala 83:49]
  wire  _dataArb_io_in_3_valid_T_45 = ((_dataArb_io_in_3_valid_res_T | (io_cpu_req_bits_cmd == 5'h11)) | _s0_read_T_3)
     | _s0_read_T_21; // @[Consts.scala 83:76]
  wire  _dataArb_io_in_3_valid_T_49 = _dataArb_io_in_3_valid_T_45 & _dataArb_io_in_3_valid_T_24; // @[DCache.scala 1086:23]
  wire  _dataArb_io_in_3_valid_T_50 = s0_read | _dataArb_io_in_3_valid_T_49; // @[DCache.scala 1085:21]
  wire  _dataArb_io_in_3_valid_T_56 = io_cpu_req_valid & res; // @[DCache.scala 212:46]
  wire  _T_4 = (~dataArb_io_in_3_ready) & s0_read; // @[DCache.scala 218:33]
  wire  _GEN_28 = _T_4 ? 1'h0 : _io_cpu_req_ready_T_4; // @[DCache.scala 218:45 DCache.scala 218:64 DCache.scala 203:20]
  wire  _s1_did_read_T_52 = dataArb_io_in_3_ready & (io_cpu_req_valid & _dataArb_io_in_3_valid_T_50); // @[DCache.scala 219:54]
  reg  s1_did_read; // @[Reg.scala 15:16]
  wire  _GEN_30 = _T ? 1'h0 : _GEN_28; // @[DCache.scala 226:34 DCache.scala 226:53]
  wire  _T_10 = ((~tlb_io_req_ready) & (~tlb_io_ptw_resp_valid)) & (~io_cpu_req_bits_phys); // @[DCache.scala 234:53]
  wire  _GEN_31 = _T_10 ? 1'h0 : _GEN_30; // @[DCache.scala 234:79 DCache.scala 234:98]
  wire [19:0] s1_paddr_right = tlb_io_resp_paddr[31:12]; // @[DCache.scala 250:99]
  wire [11:0] s1_paddr_left = s1_req_addr[11:0]; // @[DCache.scala 250:125]
  wire [31:0] s1_paddr = {s1_paddr_right,s1_paddr_left}; // @[Cat.scala 29:58]
  wire [1:0] s1_victim_way_x32 = lfsr[1:0]; // @[package.scala 143:13]
  wire  _T_19 = metaArb_io_out_valid & metaArb_io_out_bits_write; // @[DCache.scala 262:27]
  wire [21:0] _s1_meta_uncorrected_WIRE = tag_array_RW0_rdata_0;
  wire [19:0] s1_meta_uncorrected_0_tag = _s1_meta_uncorrected_WIRE[19:0]; // @[DCache.scala 267:80]
  wire [1:0] s1_meta_uncorrected_0_coh_state = _s1_meta_uncorrected_WIRE[21:20]; // @[DCache.scala 267:80]
  wire [21:0] _s1_meta_uncorrected_WIRE_1 = tag_array_RW0_rdata_1;
  wire [19:0] s1_meta_uncorrected_1_tag = _s1_meta_uncorrected_WIRE_1[19:0]; // @[DCache.scala 267:80]
  wire [1:0] s1_meta_uncorrected_1_coh_state = _s1_meta_uncorrected_WIRE_1[21:20]; // @[DCache.scala 267:80]
  wire [21:0] _s1_meta_uncorrected_WIRE_2 = tag_array_RW0_rdata_2;
  wire [19:0] s1_meta_uncorrected_2_tag = _s1_meta_uncorrected_WIRE_2[19:0]; // @[DCache.scala 267:80]
  wire [1:0] s1_meta_uncorrected_2_coh_state = _s1_meta_uncorrected_WIRE_2[21:20]; // @[DCache.scala 267:80]
  wire [21:0] _s1_meta_uncorrected_WIRE_3 = tag_array_RW0_rdata_3;
  wire [19:0] s1_meta_uncorrected_3_tag = _s1_meta_uncorrected_WIRE_3[19:0]; // @[DCache.scala 267:80]
  wire [1:0] s1_meta_uncorrected_3_coh_state = _s1_meta_uncorrected_WIRE_3[21:20]; // @[DCache.scala 267:80]
  wire [19:0] s1_tag = s1_paddr[31:12]; // @[DCache.scala 268:29]
  wire  _s1_meta_hit_way_T = s1_meta_uncorrected_0_coh_state > 2'h0; // @[Metadata.scala 50:45]
  wire  _s1_meta_hit_way_T_1 = s1_meta_uncorrected_0_tag == s1_tag; // @[DCache.scala 269:83]
  wire  s1_meta_hit_way_left_left = _s1_meta_hit_way_T & (s1_meta_uncorrected_0_tag == s1_tag); // @[DCache.scala 269:74]
  wire  _s1_meta_hit_way_T_2 = s1_meta_uncorrected_1_coh_state > 2'h0; // @[Metadata.scala 50:45]
  wire  _s1_meta_hit_way_T_3 = s1_meta_uncorrected_1_tag == s1_tag; // @[DCache.scala 269:83]
  wire  s1_meta_hit_way_left_right = _s1_meta_hit_way_T_2 & (s1_meta_uncorrected_1_tag == s1_tag); // @[DCache.scala 269:74]
  wire  _s1_meta_hit_way_T_4 = s1_meta_uncorrected_2_coh_state > 2'h0; // @[Metadata.scala 50:45]
  wire  _s1_meta_hit_way_T_5 = s1_meta_uncorrected_2_tag == s1_tag; // @[DCache.scala 269:83]
  wire  s1_meta_hit_way_right_left = _s1_meta_hit_way_T_4 & (s1_meta_uncorrected_2_tag == s1_tag); // @[DCache.scala 269:74]
  wire  _s1_meta_hit_way_T_6 = s1_meta_uncorrected_3_coh_state > 2'h0; // @[Metadata.scala 50:45]
  wire  _s1_meta_hit_way_T_7 = s1_meta_uncorrected_3_tag == s1_tag; // @[DCache.scala 269:83]
  wire  s1_meta_hit_way_right_right = _s1_meta_hit_way_T_6 & (s1_meta_uncorrected_3_tag == s1_tag); // @[DCache.scala 269:74]
  wire [3:0] s1_meta_hit_way = {s1_meta_hit_way_right_right,s1_meta_hit_way_right_left,s1_meta_hit_way_left_right,
    s1_meta_hit_way_left_left}; // @[Cat.scala 29:58]
  wire [1:0] _s1_meta_hit_state_T_3 = _s1_meta_hit_way_T_1 ? s1_meta_uncorrected_0_coh_state : 2'h0; // @[DCache.scala 271:41]
  wire [1:0] _s1_meta_hit_state_T_7 = _s1_meta_hit_way_T_3 ? s1_meta_uncorrected_1_coh_state : 2'h0; // @[DCache.scala 271:41]
  wire [1:0] _s1_meta_hit_state_T_11 = _s1_meta_hit_way_T_5 ? s1_meta_uncorrected_2_coh_state : 2'h0; // @[DCache.scala 271:41]
  wire [1:0] _s1_meta_hit_state_T_15 = _s1_meta_hit_way_T_7 ? s1_meta_uncorrected_3_coh_state : 2'h0; // @[DCache.scala 271:41]
  wire [1:0] _s1_meta_hit_state_T_16 = _s1_meta_hit_state_T_3 | _s1_meta_hit_state_T_7; // @[DCache.scala 272:19]
  wire [1:0] _s1_meta_hit_state_T_17 = _s1_meta_hit_state_T_16 | _s1_meta_hit_state_T_11; // @[DCache.scala 272:19]
  wire [1:0] s1_meta_hit_state_state = _s1_meta_hit_state_T_17 | _s1_meta_hit_state_T_15; // @[DCache.scala 272:19]
  wire  s2_hit_valid = s2_hit_state_state > 2'h0; // @[Metadata.scala 50:45]
  reg [3:0] s2_hit_way; // @[Reg.scala 15:16]
  reg [1:0] s2_victim_way_r; // @[Reg.scala 15:16]
  wire [3:0] _s2_victim_way_T_1 = 4'h1 << s2_victim_way_r; // @[OneHot.scala 58:35]
  wire [3:0] s2_victim_way = s2_hit_valid ? s2_hit_way : _s2_victim_way_T_1; // @[DCache.scala 383:26]
  reg [3:0] s2_probe_way; // @[Reg.scala 15:16]
  wire [3:0] releaseWay = _T_275 ? s2_victim_way : s2_probe_way; // @[DCache.scala 783:81 DCache.scala 790:18 DCache.scala 735:14]
  wire [3:0] s1_data_way_x34 = inWriteback ? releaseWay : s1_meta_hit_way; // @[DCache.scala 275:61]
  wire [7:0] tl_d_data_encoded_left_left_left = auto_out_d_bits_data[7:0]; // @[package.scala 183:50]
  wire [7:0] tl_d_data_encoded_left_left_right = auto_out_d_bits_data[15:8]; // @[package.scala 183:50]
  wire [7:0] tl_d_data_encoded_left_right_left = auto_out_d_bits_data[23:16]; // @[package.scala 183:50]
  wire [7:0] tl_d_data_encoded_left_right_right = auto_out_d_bits_data[31:24]; // @[package.scala 183:50]
  wire [7:0] tl_d_data_encoded_right_left_left = auto_out_d_bits_data[39:32]; // @[package.scala 183:50]
  wire [7:0] tl_d_data_encoded_right_left_right = auto_out_d_bits_data[47:40]; // @[package.scala 183:50]
  wire [7:0] tl_d_data_encoded_right_right_left = auto_out_d_bits_data[55:48]; // @[package.scala 183:50]
  wire [7:0] tl_d_data_encoded_right_right_right = auto_out_d_bits_data[63:56]; // @[package.scala 183:50]
  wire [31:0] tl_d_data_encoded_left = {tl_d_data_encoded_left_right_right,tl_d_data_encoded_left_right_left,
    tl_d_data_encoded_left_left_right,tl_d_data_encoded_left_left_left}; // @[Cat.scala 29:58]
  wire [31:0] tl_d_data_encoded_right = {tl_d_data_encoded_right_right_right,tl_d_data_encoded_right_right_left,
    tl_d_data_encoded_right_left_right,tl_d_data_encoded_right_left_left}; // @[Cat.scala 29:58]
  wire [63:0] _tl_d_data_encoded_T = {tl_d_data_encoded_right_right_right,tl_d_data_encoded_right_right_left,
    tl_d_data_encoded_right_left_right,tl_d_data_encoded_right_left_left,tl_d_data_encoded_left_right_right,
    tl_d_data_encoded_left_right_left,tl_d_data_encoded_left_left_right,tl_d_data_encoded_left_left_left}; // @[Cat.scala 29:58]
  wire [7:0] _T_28 = ~io_cpu_s1_data_mask; // @[DCache.scala 281:71]
  wire [7:0] _T_29 = s1_mask_xwr | _T_28; // @[DCache.scala 281:69]
  wire  s2_valid_x36 = s1_valid_masked & (~s1_sfence); // @[DCache.scala 283:43]
  reg [39:0] s2_req_addr; // @[DCache.scala 291:19]
  reg [6:0] s2_req_tag; // @[DCache.scala 291:19]
  reg [1:0] s2_req_size; // @[DCache.scala 291:19]
  reg  s2_req_signed; // @[DCache.scala 291:19]
  reg [1:0] s2_req_dprv; // @[DCache.scala 291:19]
  wire  _s2_cmd_flush_all_T = s2_req_cmd == 5'h5; // @[DCache.scala 292:37]
  wire  s2_cmd_flush_line = _s2_cmd_flush_all_T & (s2_req_size[0]); // @[DCache.scala 293:54]
  reg  s2_tlb_xcpt_pf_ld; // @[DCache.scala 294:24]
  reg  s2_tlb_xcpt_pf_st; // @[DCache.scala 294:24]
  reg  s2_tlb_xcpt_ae_ld; // @[DCache.scala 294:24]
  reg  s2_tlb_xcpt_ae_st; // @[DCache.scala 294:24]
  reg  s2_tlb_xcpt_ma_ld; // @[DCache.scala 294:24]
  reg  s2_tlb_xcpt_ma_st; // @[DCache.scala 294:24]
  reg  s2_pma_cacheable; // @[DCache.scala 295:19]
  reg [39:0] s2_uncached_resp_addr; // @[DCache.scala 296:34]
  wire [39:0] _GEN_57 = s1_valid_not_nacked ? {{8'd0}, s1_paddr} : s2_req_addr; // @[DCache.scala 297:48 DCache.scala 299:17 DCache.scala 291:19]
  wire [6:0] _GEN_58 = s1_valid_not_nacked ? s1_req_tag : s2_req_tag; // @[DCache.scala 297:48 DCache.scala 298:12 DCache.scala 291:19]
  wire [4:0] _GEN_59 = s1_valid_not_nacked ? s1_req_cmd : s2_req_cmd; // @[DCache.scala 297:48 DCache.scala 298:12 DCache.scala 291:19]
  wire [1:0] _GEN_60 = s1_valid_not_nacked ? s1_req_size : s2_req_size; // @[DCache.scala 297:48 DCache.scala 298:12 DCache.scala 291:19]
  wire  _GEN_61 = s1_valid_not_nacked ? s1_req_signed : s2_req_signed; // @[DCache.scala 297:48 DCache.scala 298:12 DCache.scala 291:19]
  reg [39:0] s2_vaddr_r; // @[Reg.scala 15:16]
  wire [27:0] s2_vaddr_right = s2_vaddr_r[39:12]; // @[DCache.scala 303:84]
  wire [11:0] s2_vaddr_left = s2_req_addr[11:0]; // @[DCache.scala 303:109]
  wire [39:0] s2_vaddr = {s2_vaddr_right,s2_vaddr_left}; // @[Cat.scala 29:58]
  wire  en = (s1_valid | inWriteback) | io_cpu_replay_next; // @[DCache.scala 318:38]
  wire  _s2_data_word_en_T_1 = ~s1_did_read ? 1'h0 : 1'h1; // @[DCache.scala 319:63]
  wire  word_en = inWriteback | _s2_data_word_en_T_1; // @[DCache.scala 319:22]
  wire [63:0] s1_all_data_ways_0 = data_io_resp_0; // @[DCache.scala 277:29 DCache.scala 277:29]
  wire [63:0] s1_all_data_ways_1 = data_io_resp_1; // @[DCache.scala 277:29 DCache.scala 277:29]
  wire [63:0] s1_all_data_ways_2 = data_io_resp_2; // @[DCache.scala 277:29 DCache.scala 277:29]
  wire [63:0] s1_all_data_ways_3 = data_io_resp_3; // @[DCache.scala 277:29 DCache.scala 277:29]
  wire  s1_word_en = ~io_cpu_replay_next ? word_en : 1'h1; // @[DCache.scala 329:27]
  wire  grantIsUncachedData = auto_out_d_bits_opcode == 3'h1; // @[package.scala 15:47]
  reg  blockUncachedGrant; // @[DCache.scala 693:33]
  wire  _T_259 = grantIsUncachedData & (blockUncachedGrant | s1_valid); // @[DCache.scala 695:31]
  wire  grantIsRefill = auto_out_d_bits_opcode == 3'h5; // @[DCache.scala 609:29]
  wire  _T_256 = ~dataArb_io_in_1_ready; // @[DCache.scala 665:26]
  wire  _T_257 = grantIsRefill & (~dataArb_io_in_1_ready); // @[DCache.scala 665:23]
  wire  _grantIsCached_T = auto_out_d_bits_opcode == 3'h4; // @[package.scala 15:47]
  wire  grantIsCached = _grantIsCached_T | grantIsRefill; // @[package.scala 64:59]
  reg [8:0] counter; // @[Edges.scala 230:27]
  wire  d_first = counter == 9'h0; // @[Edges.scala 232:25]
  wire  canAcceptCachedGrant = ~_T_275; // @[DCache.scala 613:30]
  wire  _tl_out_d_ready_T_3 = grantIsCached ? ((~d_first) | auto_out_e_ready) & canAcceptCachedGrant : 1'h1; // @[DCache.scala 614:24]
  wire  _GEN_232 = _T_257 ? 1'h0 : _tl_out_d_ready_T_3; // @[DCache.scala 665:51 DCache.scala 667:20 DCache.scala 614:18]
  wire  tl_out__d_ready = _T_259 ? 1'h0 : _GEN_232; // @[DCache.scala 695:68 DCache.scala 696:22]
  wire  _T_236 = tl_out__d_ready & auto_out_d_valid; // @[Decoupled.scala 40:37]
  wire  _T_232 = auto_out_d_bits_opcode == 3'h0; // @[package.scala 15:47]
  wire  _T_233 = auto_out_d_bits_opcode == 3'h2; // @[package.scala 15:47]
  wire  grantIsUncached = (grantIsUncachedData | _T_232) | _T_233; // @[package.scala 64:59]
  wire [4:0] _GEN_188 = grantIsUncachedData ? 5'h10 : {{1'd0}, s1_data_way_x34}; // @[DCache.scala 634:34 DCache.scala 637:25]
  wire [4:0] _GEN_197 = grantIsUncached ? _GEN_188 : {{1'd0}, s1_data_way_x34}; // @[DCache.scala 627:35]
  wire [4:0] _GEN_210 = grantIsCached ? {{1'd0}, s1_data_way_x34} : _GEN_197; // @[DCache.scala 618:26]
  wire [4:0] s1_data_way = _T_236 ? _GEN_210 : {{1'd0}, s1_data_way_x34}; // @[DCache.scala 617:26]
  wire [4:0] _s2_data_T_1 = s1_word_en ? s1_data_way : 5'h0; // @[DCache.scala 331:28]
  wire [63:0] _s2_data_T_7 = _s2_data_T_1[0] ? s1_all_data_ways_0 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _s2_data_T_8 = _s2_data_T_1[1] ? s1_all_data_ways_1 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _s2_data_T_9 = _s2_data_T_1[2] ? s1_all_data_ways_2 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _s2_data_T_10 = _s2_data_T_1[3] ? s1_all_data_ways_3 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _s2_data_T_11 = _s2_data_T_1[4] ? _tl_d_data_encoded_T : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _s2_data_T_12 = _s2_data_T_7 | _s2_data_T_8; // @[Mux.scala 27:72]
  wire [63:0] _s2_data_T_13 = _s2_data_T_12 | _s2_data_T_9; // @[Mux.scala 27:72]
  wire [63:0] _s2_data_T_14 = _s2_data_T_13 | _s2_data_T_10; // @[Mux.scala 27:72]
  wire [63:0] _s2_data_T_15 = _s2_data_T_14 | _s2_data_T_11; // @[Mux.scala 27:72]
  reg [63:0] s2_data; // @[Reg.scala 15:16]
  wire [7:0] s2_data_uncorrected_left_left_left = s2_data[7:0]; // @[package.scala 183:50]
  wire [7:0] s2_data_uncorrected_left_left_right = s2_data[15:8]; // @[package.scala 183:50]
  wire [7:0] s2_data_uncorrected_left_right_left = s2_data[23:16]; // @[package.scala 183:50]
  wire [7:0] s2_data_uncorrected_left_right_right = s2_data[31:24]; // @[package.scala 183:50]
  wire [7:0] s2_data_uncorrected_right_left_left = s2_data[39:32]; // @[package.scala 183:50]
  wire [7:0] s2_data_uncorrected_right_left_right = s2_data[47:40]; // @[package.scala 183:50]
  wire [7:0] s2_data_uncorrected_right_right_left = s2_data[55:48]; // @[package.scala 183:50]
  wire [7:0] s2_data_uncorrected_right_right_right = s2_data[63:56]; // @[package.scala 183:50]
  wire [31:0] s2_data_corrected_left = {s2_data_uncorrected_left_right_right,s2_data_uncorrected_left_right_left,
    s2_data_uncorrected_left_left_right,s2_data_uncorrected_left_left_left}; // @[Cat.scala 29:58]
  wire [31:0] s2_data_corrected_right = {s2_data_uncorrected_right_right_right,s2_data_uncorrected_right_right_left,
    s2_data_uncorrected_right_left_right,s2_data_uncorrected_right_left_left}; // @[Cat.scala 29:58]
  wire [63:0] s2_data_corrected = {s2_data_uncorrected_right_right_right,s2_data_uncorrected_right_right_left,
    s2_data_uncorrected_right_left_right,s2_data_uncorrected_right_left_left,s2_data_uncorrected_left_right_right,
    s2_data_uncorrected_left_right_left,s2_data_uncorrected_left_left_right,s2_data_uncorrected_left_left_left}; // @[Cat.scala 29:58]
  wire  s2_valid_flush_line = s2_valid_hit_maybe_flush_pre_data_ecc_and_waw & s2_cmd_flush_line; // @[DCache.scala 371:75]
  wire  s2_valid_miss = (s2_valid_masked & s2_readwrite) & (~s2_hit); // @[DCache.scala 375:73]
  wire  s2_uncached = ~s2_pma_cacheable; // @[DCache.scala 376:21]
  wire  _s2_valid_cached_miss_T = ~s2_uncached; // @[DCache.scala 377:47]
  wire  _s2_valid_cached_miss_T_2 = |uncachedInFlight_0; // @[DCache.scala 377:88]
  wire  s2_valid_cached_miss = (s2_valid_miss & (~s2_uncached)) & (~(|uncachedInFlight_0)); // @[DCache.scala 377:60]
  wire  s2_want_victimize = s2_valid_cached_miss | s2_valid_flush_line; // @[DCache.scala 379:79]
  wire  s2_valid_uncached_pending = (s2_valid_miss & s2_uncached) & (~(&uncachedInFlight_0)); // @[DCache.scala 382:64]
  reg [19:0] s2_victim_tag_r; // @[Reg.scala 15:16]
  wire [19:0] s2_victim_tag = s2_valid_flush_line ? s2_req_addr[31:12] : s2_victim_tag_r; // @[DCache.scala 384:26]
  reg [1:0] s2_victim_state_r_state; // @[Reg.scala 15:16]
  wire [1:0] s2_victim_state_state = s2_hit_valid ? s2_hit_state_state : s2_victim_state_r_state; // @[DCache.scala 385:28]
  wire [2:0] _T_98 = _T_96 ? 3'h5 : 3'h0; // @[Misc.scala 37:36]
  wire [2:0] _T_102 = _T_100 ? 3'h2 : _T_98; // @[Misc.scala 37:36]
  wire [2:0] _T_106 = _T_104 ? 3'h1 : _T_102; // @[Misc.scala 37:36]
  wire [2:0] _T_110 = _T_108 ? 3'h1 : _T_106; // @[Misc.scala 37:36]
  wire [2:0] _T_114 = _T_112 ? 3'h5 : _T_110; // @[Misc.scala 37:36]
  wire [2:0] _T_118 = _T_116 ? 3'h4 : _T_114; // @[Misc.scala 37:36]
  wire [1:0] _T_119 = _T_116 ? 2'h1 : 2'h0; // @[Misc.scala 37:63]
  wire [2:0] _T_122 = _T_120 ? 3'h0 : _T_118; // @[Misc.scala 37:36]
  wire [1:0] _T_123 = _T_120 ? 2'h1 : _T_119; // @[Misc.scala 37:63]
  wire [2:0] _T_126 = _T_124 ? 3'h0 : _T_122; // @[Misc.scala 37:36]
  wire [1:0] _T_127 = _T_124 ? 2'h1 : _T_123; // @[Misc.scala 37:63]
  wire [2:0] _T_130 = _T_128 ? 3'h5 : _T_126; // @[Misc.scala 37:36]
  wire [1:0] _T_131 = _T_128 ? 2'h0 : _T_127; // @[Misc.scala 37:63]
  wire [2:0] _T_134 = _T_132 ? 3'h4 : _T_130; // @[Misc.scala 37:36]
  wire [1:0] _T_135 = _T_132 ? 2'h1 : _T_131; // @[Misc.scala 37:63]
  wire [2:0] _T_138 = _T_136 ? 3'h3 : _T_134; // @[Misc.scala 37:36]
  wire [1:0] _T_139 = _T_136 ? 2'h2 : _T_135; // @[Misc.scala 37:63]
  wire [2:0] s2_report_param = _T_140 ? 3'h3 : _T_138; // @[Misc.scala 37:36]
  wire [1:0] probeNewCoh_state = _T_140 ? 2'h2 : _T_139; // @[Misc.scala 37:63]
  wire [3:0] _T_147 = {2'h2,s2_victim_state_state}; // @[Cat.scala 29:58]
  wire  _T_160 = 4'h8 == _T_147; // @[Misc.scala 55:20]
  wire [2:0] _T_162 = _T_160 ? 3'h5 : 3'h0; // @[Misc.scala 37:36]
  wire  _T_164 = 4'h9 == _T_147; // @[Misc.scala 55:20]
  wire [2:0] _T_166 = _T_164 ? 3'h2 : _T_162; // @[Misc.scala 37:36]
  wire  _T_168 = 4'ha == _T_147; // @[Misc.scala 55:20]
  wire [2:0] _T_170 = _T_168 ? 3'h1 : _T_166; // @[Misc.scala 37:36]
  wire  _T_172 = 4'hb == _T_147; // @[Misc.scala 55:20]
  wire [2:0] _T_174 = _T_172 ? 3'h1 : _T_170; // @[Misc.scala 37:36]
  wire  _T_176 = 4'h4 == _T_147; // @[Misc.scala 55:20]
  wire  _T_177 = _T_176 ? 1'h0 : _T_172; // @[Misc.scala 37:9]
  wire [2:0] _T_178 = _T_176 ? 3'h5 : _T_174; // @[Misc.scala 37:36]
  wire  _T_180 = 4'h5 == _T_147; // @[Misc.scala 55:20]
  wire  _T_181 = _T_180 ? 1'h0 : _T_177; // @[Misc.scala 37:9]
  wire [2:0] _T_182 = _T_180 ? 3'h4 : _T_178; // @[Misc.scala 37:36]
  wire [1:0] _T_183 = _T_180 ? 2'h1 : 2'h0; // @[Misc.scala 37:63]
  wire  _T_184 = 4'h6 == _T_147; // @[Misc.scala 55:20]
  wire  _T_185 = _T_184 ? 1'h0 : _T_181; // @[Misc.scala 37:9]
  wire [2:0] _T_186 = _T_184 ? 3'h0 : _T_182; // @[Misc.scala 37:36]
  wire [1:0] _T_187 = _T_184 ? 2'h1 : _T_183; // @[Misc.scala 37:63]
  wire  _T_188 = 4'h7 == _T_147; // @[Misc.scala 55:20]
  wire [2:0] _T_190 = _T_188 ? 3'h0 : _T_186; // @[Misc.scala 37:36]
  wire [1:0] _T_191 = _T_188 ? 2'h1 : _T_187; // @[Misc.scala 37:63]
  wire  _T_192 = 4'h0 == _T_147; // @[Misc.scala 55:20]
  wire  _T_193 = _T_192 ? 1'h0 : _T_188 | _T_185; // @[Misc.scala 37:9]
  wire [2:0] _T_194 = _T_192 ? 3'h5 : _T_190; // @[Misc.scala 37:36]
  wire [1:0] _T_195 = _T_192 ? 2'h0 : _T_191; // @[Misc.scala 37:63]
  wire  _T_196 = 4'h1 == _T_147; // @[Misc.scala 55:20]
  wire  _T_197 = _T_196 ? 1'h0 : _T_193; // @[Misc.scala 37:9]
  wire [2:0] _T_198 = _T_196 ? 3'h4 : _T_194; // @[Misc.scala 37:36]
  wire [1:0] _T_199 = _T_196 ? 2'h1 : _T_195; // @[Misc.scala 37:63]
  wire  _T_200 = 4'h2 == _T_147; // @[Misc.scala 55:20]
  wire  _T_201 = _T_200 ? 1'h0 : _T_197; // @[Misc.scala 37:9]
  wire [2:0] _T_202 = _T_200 ? 3'h3 : _T_198; // @[Misc.scala 37:36]
  wire [1:0] _T_203 = _T_200 ? 2'h2 : _T_199; // @[Misc.scala 37:63]
  wire  _T_204 = 4'h3 == _T_147; // @[Misc.scala 55:20]
  wire  s2_victim_dirty = _T_204 | _T_201; // @[Misc.scala 37:9]
  wire [2:0] s2_shrink_param = _T_204 ? 3'h3 : _T_202; // @[Misc.scala 37:36]
  wire [1:0] voluntaryNewCoh_state = _T_204 ? 2'h2 : _T_203; // @[Misc.scala 37:63]
  wire  s2_dont_nack_uncached = s2_valid_uncached_pending & auto_out_a_ready; // @[DCache.scala 391:57]
  wire  _s2_dont_nack_misc_T_10 = s2_req_cmd == 5'h17; // @[DCache.scala 395:17]
  wire  s2_dont_nack_misc = s2_valid_masked & _s2_dont_nack_misc_T_10; // @[DCache.scala 392:61]
  wire  _io_cpu_s2_nack_T_4 = ~s2_valid_hit_pre_data_ecc_and_waw; // @[DCache.scala 396:89]
  wire [27:0] metaArb_io_in_1_bits_addr_right = io_cpu_req_bits_addr[39:12]; // @[DCache.scala 405:58]
  wire [11:0] metaArb_io_in_2_bits_addr_left = s2_vaddr[11:0]; // @[DCache.scala 417:80]
  wire [19:0] metaArb_io_in_2_bits_data_meta_tag = s2_req_addr[31:12]; // @[HellaCache.scala 282:20 HellaCache.scala 283:14]
  wire  _lrscBackingOff_T = lrscCount > 7'h0; // @[DCache.scala 425:34]
  wire  lrscBackingOff = (lrscCount > 7'h0) & (~lrscValid); // @[DCache.scala 425:38]
  reg [33:0] lrscAddr; // @[DCache.scala 426:21]
  wire  lrscAddrMatch = lrscAddr == (s2_req_addr[39:6]); // @[DCache.scala 427:32]
  wire  s2_sc_fail = _s2_write_T_3 & (~(lrscValid & lrscAddrMatch)); // @[DCache.scala 428:26]
  wire  _T_211 = ((s2_valid_hit_pre_data_ecc_and_waw & _c_cat_T_47) & _io_cpu_req_ready_T_1) | s2_valid_cached_miss; // @[DCache.scala 429:54]
  wire [6:0] _lrscCount_T = s2_hit ? 7'h4f : 7'h0; // @[DCache.scala 430:21]
  wire [6:0] _GEN_120 = _T_211 ? _lrscCount_T : lrscCount; // @[DCache.scala 429:99 DCache.scala 430:15 DCache.scala 423:22]
  wire [6:0] _lrscCount_T_2 = lrscCount - 7'h1; // @[DCache.scala 433:49]
  wire  _T_215 = s2_valid_masked & lrscValid; // @[DCache.scala 434:29]
  wire  _pstore1_cmd_T = s1_valid_not_nacked & s1_write; // @[DCache.scala 443:63]
  reg [4:0] pstore1_cmd; // @[Reg.scala 15:16]
  reg [63:0] pstore1_data; // @[Reg.scala 15:16]
  reg [3:0] pstore1_way; // @[Reg.scala 15:16]
  wire  _pstore1_rmw_T_49 = s1_write & _s1_write_T_1; // @[DCache.scala 1086:23]
  wire  _pstore1_rmw_T_50 = s1_read | _pstore1_rmw_T_49; // @[DCache.scala 1085:21]
  reg  pstore1_rmw_r; // @[Reg.scala 15:16]
  wire  _pstore1_merge_T = s2_valid_hit_pre_data_ecc_and_waw & s2_write; // @[DCache.scala 441:46]
  wire  _pstore1_merge_T_2 = (s2_valid_hit_pre_data_ecc_and_waw & s2_write) & (~s2_sc_fail); // @[DCache.scala 441:58]
  wire  pstore_drain_opportunistic = ~_dataArb_io_in_3_valid_T_56; // @[DCache.scala 453:36]
  reg  pstore_drain_on_miss_REG; // @[DCache.scala 454:56]
  wire  pstore_drain_on_miss = releaseInFlight | pstore_drain_on_miss_REG; // @[DCache.scala 454:46]
  wire  pstore1_valid = _pstore1_merge_T_2 | pstore1_held; // @[DCache.scala 458:38]
  wire  pstore_drain_structural = (pstore1_valid_likely & pstore2_valid) & ((s1_valid & s1_write) | pstore1_rmw_r); // @[DCache.scala 460:71]
  wire  _T_219 = _pstore1_merge_T | pstore1_held; // @[DCache.scala 457:96]
  wire  _pstore_drain_T_10 = ((_T_219 & (~pstore1_rmw_r)) | pstore2_valid) & (pstore_drain_opportunistic |
    pstore_drain_on_miss); // @[DCache.scala 469:76]
  wire  pstore_drain = pstore_drain_structural | _pstore_drain_T_10; // @[DCache.scala 468:48]
  wire  _pstore1_held_T_9 = ~pstore_drain; // @[DCache.scala 472:91]
  wire  advance_pstore1 = pstore1_valid & (pstore2_valid == pstore_drain); // @[DCache.scala 473:61]
  reg [3:0] pstore2_way; // @[Reg.scala 15:16]
  wire [63:0] pstore1_storegen_data = amoalu_io_out;
  reg [7:0] pstore2_storegen_data_left_left_left; // @[Reg.scala 15:16]
  reg [7:0] pstore2_storegen_data_left_left_right; // @[Reg.scala 15:16]
  reg [7:0] pstore2_storegen_data_left_right_left; // @[Reg.scala 15:16]
  reg [7:0] pstore2_storegen_data_left_right_right; // @[Reg.scala 15:16]
  reg [7:0] pstore2_storegen_data_right_left_left; // @[Reg.scala 15:16]
  reg [7:0] pstore2_storegen_data_right_left_right; // @[Reg.scala 15:16]
  reg [7:0] pstore2_storegen_data_right_right_left; // @[Reg.scala 15:16]
  reg [7:0] pstore2_storegen_data_right_right_right; // @[Reg.scala 15:16]
  wire [63:0] pstore2_storegen_data = {pstore2_storegen_data_right_right_right,pstore2_storegen_data_right_right_left,
    pstore2_storegen_data_right_left_right,pstore2_storegen_data_right_left_left,pstore2_storegen_data_left_right_right,
    pstore2_storegen_data_left_right_left,pstore2_storegen_data_left_left_right,pstore2_storegen_data_left_left_left}; // @[Cat.scala 29:58]
  wire [7:0] _pstore2_storegen_mask_mask_T = ~pstore1_mask; // @[DCache.scala 485:37]
  wire [7:0] _pstore2_storegen_mask_mask_T_2 = ~_pstore2_storegen_mask_mask_T; // @[DCache.scala 485:15]
  wire [39:0] _dataArb_io_in_0_bits_addr_T = pstore2_valid ? pstore2_addr : pstore1_addr; // @[DCache.scala 500:36]
  wire [63:0] _dataArb_io_in_0_bits_wdata_T = pstore2_valid ? pstore2_storegen_data : pstore1_data; // @[DCache.scala 502:63]
  wire [7:0] dataArb_io_in_0_bits_wdata_left_left_left = _dataArb_io_in_0_bits_wdata_T[7:0]; // @[package.scala 183:50]
  wire [7:0] dataArb_io_in_0_bits_wdata_left_left_right = _dataArb_io_in_0_bits_wdata_T[15:8]; // @[package.scala 183:50]
  wire [7:0] dataArb_io_in_0_bits_wdata_left_right_left = _dataArb_io_in_0_bits_wdata_T[23:16]; // @[package.scala 183:50]
  wire [7:0] dataArb_io_in_0_bits_wdata_left_right_right = _dataArb_io_in_0_bits_wdata_T[31:24]; // @[package.scala 183:50]
  wire [7:0] dataArb_io_in_0_bits_wdata_right_left_left = _dataArb_io_in_0_bits_wdata_T[39:32]; // @[package.scala 183:50]
  wire [7:0] dataArb_io_in_0_bits_wdata_right_left_right = _dataArb_io_in_0_bits_wdata_T[47:40]; // @[package.scala 183:50]
  wire [7:0] dataArb_io_in_0_bits_wdata_right_right_left = _dataArb_io_in_0_bits_wdata_T[55:48]; // @[package.scala 183:50]
  wire [7:0] dataArb_io_in_0_bits_wdata_right_right_right = _dataArb_io_in_0_bits_wdata_T[63:56]; // @[package.scala 183:50]
  wire [31:0] dataArb_io_in_0_bits_wdata_left = {dataArb_io_in_0_bits_wdata_left_right_right,
    dataArb_io_in_0_bits_wdata_left_right_left,dataArb_io_in_0_bits_wdata_left_left_right,
    dataArb_io_in_0_bits_wdata_left_left_left}; // @[Cat.scala 29:58]
  wire [31:0] dataArb_io_in_0_bits_wdata_right = {dataArb_io_in_0_bits_wdata_right_right_right,
    dataArb_io_in_0_bits_wdata_right_right_left,dataArb_io_in_0_bits_wdata_right_left_right,
    dataArb_io_in_0_bits_wdata_right_left_left}; // @[Cat.scala 29:58]
  wire [7:0] _dataArb_io_in_0_bits_eccMask_T = pstore2_valid ? mask : pstore1_mask; // @[DCache.scala 504:47]
  wire  dataArb_io_in_0_bits_eccMask_left_left_left = |(_dataArb_io_in_0_bits_eccMask_T[0]); // @[DCache.scala 1076:66]
  wire  dataArb_io_in_0_bits_eccMask_left_left_right = |(_dataArb_io_in_0_bits_eccMask_T[1]); // @[DCache.scala 1076:66]
  wire  dataArb_io_in_0_bits_eccMask_left_right_left = |(_dataArb_io_in_0_bits_eccMask_T[2]); // @[DCache.scala 1076:66]
  wire  dataArb_io_in_0_bits_eccMask_left_right_right = |(_dataArb_io_in_0_bits_eccMask_T[3]); // @[DCache.scala 1076:66]
  wire  dataArb_io_in_0_bits_eccMask_right_left_left = |(_dataArb_io_in_0_bits_eccMask_T[4]); // @[DCache.scala 1076:66]
  wire  dataArb_io_in_0_bits_eccMask_right_left_right = |(_dataArb_io_in_0_bits_eccMask_T[5]); // @[DCache.scala 1076:66]
  wire  dataArb_io_in_0_bits_eccMask_right_right_left = |(_dataArb_io_in_0_bits_eccMask_T[6]); // @[DCache.scala 1076:66]
  wire  dataArb_io_in_0_bits_eccMask_right_right_right = |(_dataArb_io_in_0_bits_eccMask_T[7]); // @[DCache.scala 1076:66]
  wire [3:0] dataArb_io_in_0_bits_eccMask_left = {dataArb_io_in_0_bits_eccMask_left_right_right,
    dataArb_io_in_0_bits_eccMask_left_right_left,dataArb_io_in_0_bits_eccMask_left_left_right,
    dataArb_io_in_0_bits_eccMask_left_left_left}; // @[Cat.scala 29:58]
  wire [3:0] dataArb_io_in_0_bits_eccMask_right = {dataArb_io_in_0_bits_eccMask_right_right_right,
    dataArb_io_in_0_bits_eccMask_right_right_left,dataArb_io_in_0_bits_eccMask_right_left_right,
    dataArb_io_in_0_bits_eccMask_right_left_left}; // @[Cat.scala 29:58]
  wire  _a_source_T = ~uncachedInFlight_0; // @[DCache.scala 524:34]
  wire [1:0] _a_source_T_1 = {_a_source_T, 1'h0}; // @[DCache.scala 524:59]
  wire  a_source = _a_source_T_1[0] ? 1'h0 : 1'h1; // @[Mux.scala 47:69]
  wire [39:0] acquire_address = {s2_req_addr[39:6], 6'h0}; // @[DCache.scala 525:49]
  wire [22:0] a_mask = {{15'd0}, pstore1_mask}; // @[DCache.scala 529:29]
  wire [2:0] _get_get_mask_sizeOH_T = {{1'd0}, s2_req_size}; // @[Misc.scala 201:34]
  wire [1:0] get_get_mask_sizeOH_shiftAmount = _get_get_mask_sizeOH_T[1:0]; // @[OneHot.scala 64:49]
  wire [3:0] _get_get_mask_sizeOH_T_1 = 4'h1 << get_get_mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12]
  wire [2:0] get_get_mask_sizeOH = (_get_get_mask_sizeOH_T_1[2:0]) | 3'h1; // @[Misc.scala 201:81]
  wire  get_get_mask_sub_acc = s2_req_size >= 2'h3; // @[Misc.scala 205:21]
  wire  get_get_mask_size = get_get_mask_sizeOH[2]; // @[Misc.scala 208:26]
  wire  get_get_mask_bit = s2_req_addr[2]; // @[Misc.scala 209:26]
  wire  get_get_mask_nbit = ~get_get_mask_bit; // @[Misc.scala 210:20]
  wire  get_get_mask_sub_acc_1 = get_get_mask_sub_acc | (get_get_mask_size & get_get_mask_nbit); // @[Misc.scala 214:29]
  wire  get_get_mask_sub_acc_2 = get_get_mask_sub_acc | (get_get_mask_size & get_get_mask_bit); // @[Misc.scala 214:29]
  wire  get_get_mask_size_1 = get_get_mask_sizeOH[1]; // @[Misc.scala 208:26]
  wire  get_get_mask_bit_1 = s2_req_addr[1]; // @[Misc.scala 209:26]
  wire  get_get_mask_nbit_1 = ~get_get_mask_bit_1; // @[Misc.scala 210:20]
  wire  get_get_mask_sub_eq_2 = get_get_mask_nbit & get_get_mask_nbit_1; // @[Misc.scala 213:27]
  wire  get_get_mask_sub_acc_3 = get_get_mask_sub_acc_1 | (get_get_mask_size_1 & get_get_mask_sub_eq_2); // @[Misc.scala 214:29]
  wire  get_get_mask_sub_eq_3 = get_get_mask_nbit & get_get_mask_bit_1; // @[Misc.scala 213:27]
  wire  get_get_mask_sub_acc_4 = get_get_mask_sub_acc_1 | (get_get_mask_size_1 & get_get_mask_sub_eq_3); // @[Misc.scala 214:29]
  wire  get_get_mask_sub_eq_4 = get_get_mask_bit & get_get_mask_nbit_1; // @[Misc.scala 213:27]
  wire  get_get_mask_sub_acc_5 = get_get_mask_sub_acc_2 | (get_get_mask_size_1 & get_get_mask_sub_eq_4); // @[Misc.scala 214:29]
  wire  get_get_mask_sub_eq_5 = get_get_mask_bit & get_get_mask_bit_1; // @[Misc.scala 213:27]
  wire  get_get_mask_sub_acc_6 = get_get_mask_sub_acc_2 | (get_get_mask_size_1 & get_get_mask_sub_eq_5); // @[Misc.scala 214:29]
  wire  get_get_mask_size_2 = get_get_mask_sizeOH[0]; // @[Misc.scala 208:26]
  wire  get_get_mask_bit_2 = s2_req_addr[0]; // @[Misc.scala 209:26]
  wire  get_get_mask_nbit_2 = ~get_get_mask_bit_2; // @[Misc.scala 210:20]
  wire  get_get_mask_eq = get_get_mask_sub_eq_2 & get_get_mask_nbit_2; // @[Misc.scala 213:27]
  wire  get_get_mask_left_left_left = get_get_mask_sub_acc_3 | (get_get_mask_size_2 & get_get_mask_eq); // @[Misc.scala 214:29]
  wire  get_get_mask_eq_1 = get_get_mask_sub_eq_2 & get_get_mask_bit_2; // @[Misc.scala 213:27]
  wire  get_get_mask_left_left_right = get_get_mask_sub_acc_3 | (get_get_mask_size_2 & get_get_mask_eq_1); // @[Misc.scala 214:29]
  wire  get_get_mask_eq_2 = get_get_mask_sub_eq_3 & get_get_mask_nbit_2; // @[Misc.scala 213:27]
  wire  get_get_mask_left_right_left = get_get_mask_sub_acc_4 | (get_get_mask_size_2 & get_get_mask_eq_2); // @[Misc.scala 214:29]
  wire  get_get_mask_eq_3 = get_get_mask_sub_eq_3 & get_get_mask_bit_2; // @[Misc.scala 213:27]
  wire  get_get_mask_left_right_right = get_get_mask_sub_acc_4 | (get_get_mask_size_2 & get_get_mask_eq_3); // @[Misc.scala 214:29]
  wire  get_get_mask_eq_4 = get_get_mask_sub_eq_4 & get_get_mask_nbit_2; // @[Misc.scala 213:27]
  wire  get_get_mask_right_left_left = get_get_mask_sub_acc_5 | (get_get_mask_size_2 & get_get_mask_eq_4); // @[Misc.scala 214:29]
  wire  get_get_mask_eq_5 = get_get_mask_sub_eq_4 & get_get_mask_bit_2; // @[Misc.scala 213:27]
  wire  get_get_mask_right_left_right = get_get_mask_sub_acc_5 | (get_get_mask_size_2 & get_get_mask_eq_5); // @[Misc.scala 214:29]
  wire  get_get_mask_eq_6 = get_get_mask_sub_eq_5 & get_get_mask_nbit_2; // @[Misc.scala 213:27]
  wire  get_get_mask_right_right_left = get_get_mask_sub_acc_6 | (get_get_mask_size_2 & get_get_mask_eq_6); // @[Misc.scala 214:29]
  wire  get_get_mask_eq_7 = get_get_mask_sub_eq_5 & get_get_mask_bit_2; // @[Misc.scala 213:27]
  wire  get_get_mask_right_right_right = get_get_mask_sub_acc_6 | (get_get_mask_size_2 & get_get_mask_eq_7); // @[Misc.scala 214:29]
  wire [7:0] get_mask = {get_get_mask_right_right_right,get_get_mask_right_right_left,get_get_mask_right_left_right,
    get_get_mask_right_left_left,get_get_mask_left_right_right,get_get_mask_left_right_left,get_get_mask_left_left_right
    ,get_get_mask_left_left_left}; // @[Cat.scala 29:58]
  wire [2:0] _atomics_T_1_opcode = 5'h4 == s2_req_cmd ? 3'h3 : 3'h0; // @[Mux.scala 80:57]
  wire [3:0] atomics_a_size = {{2'd0}, s2_req_size}; // @[Edges.scala 515:17 Edges.scala 518:15]
  wire [3:0] _atomics_T_1_size = 5'h4 == s2_req_cmd ? atomics_a_size : 4'h0; // @[Mux.scala 80:57]
  wire [31:0] atomics_a_address = s2_req_addr[31:0]; // @[Edges.scala 515:17 Edges.scala 520:15]
  wire [31:0] _atomics_T_1_address = 5'h4 == s2_req_cmd ? atomics_a_address : 32'h0; // @[Mux.scala 80:57]
  wire [7:0] _atomics_T_1_mask = 5'h4 == s2_req_cmd ? get_mask : 8'h0; // @[Mux.scala 80:57]
  wire [63:0] _atomics_T_1_data = 5'h4 == s2_req_cmd ? pstore1_data : 64'h0; // @[Mux.scala 80:57]
  wire [2:0] _atomics_T_3_opcode = 5'h9 == s2_req_cmd ? 3'h3 : _atomics_T_1_opcode; // @[Mux.scala 80:57]
  wire [2:0] _atomics_T_3_param = 5'h9 == s2_req_cmd ? 3'h0 : _atomics_T_1_opcode; // @[Mux.scala 80:57]
  wire [3:0] _atomics_T_3_size = 5'h9 == s2_req_cmd ? atomics_a_size : _atomics_T_1_size; // @[Mux.scala 80:57]
  wire  _atomics_T_3_source = 5'h9 == s2_req_cmd ? a_source : (5'h4 == s2_req_cmd) & a_source; // @[Mux.scala 80:57]
  wire [31:0] _atomics_T_3_address = 5'h9 == s2_req_cmd ? atomics_a_address : _atomics_T_1_address; // @[Mux.scala 80:57]
  wire [7:0] _atomics_T_3_mask = 5'h9 == s2_req_cmd ? get_mask : _atomics_T_1_mask; // @[Mux.scala 80:57]
  wire [63:0] _atomics_T_3_data = 5'h9 == s2_req_cmd ? pstore1_data : _atomics_T_1_data; // @[Mux.scala 80:57]
  wire [2:0] _atomics_T_5_opcode = 5'ha == s2_req_cmd ? 3'h3 : _atomics_T_3_opcode; // @[Mux.scala 80:57]
  wire [2:0] _atomics_T_5_param = 5'ha == s2_req_cmd ? 3'h1 : _atomics_T_3_param; // @[Mux.scala 80:57]
  wire [3:0] _atomics_T_5_size = 5'ha == s2_req_cmd ? atomics_a_size : _atomics_T_3_size; // @[Mux.scala 80:57]
  wire  _atomics_T_5_source = 5'ha == s2_req_cmd ? a_source : _atomics_T_3_source; // @[Mux.scala 80:57]
  wire [31:0] _atomics_T_5_address = 5'ha == s2_req_cmd ? atomics_a_address : _atomics_T_3_address; // @[Mux.scala 80:57]
  wire [7:0] _atomics_T_5_mask = 5'ha == s2_req_cmd ? get_mask : _atomics_T_3_mask; // @[Mux.scala 80:57]
  wire [63:0] _atomics_T_5_data = 5'ha == s2_req_cmd ? pstore1_data : _atomics_T_3_data; // @[Mux.scala 80:57]
  wire [2:0] _atomics_T_7_opcode = 5'hb == s2_req_cmd ? 3'h3 : _atomics_T_5_opcode; // @[Mux.scala 80:57]
  wire [2:0] _atomics_T_7_param = 5'hb == s2_req_cmd ? 3'h2 : _atomics_T_5_param; // @[Mux.scala 80:57]
  wire [3:0] _atomics_T_7_size = 5'hb == s2_req_cmd ? atomics_a_size : _atomics_T_5_size; // @[Mux.scala 80:57]
  wire  _atomics_T_7_source = 5'hb == s2_req_cmd ? a_source : _atomics_T_5_source; // @[Mux.scala 80:57]
  wire [31:0] _atomics_T_7_address = 5'hb == s2_req_cmd ? atomics_a_address : _atomics_T_5_address; // @[Mux.scala 80:57]
  wire [7:0] _atomics_T_7_mask = 5'hb == s2_req_cmd ? get_mask : _atomics_T_5_mask; // @[Mux.scala 80:57]
  wire [63:0] _atomics_T_7_data = 5'hb == s2_req_cmd ? pstore1_data : _atomics_T_5_data; // @[Mux.scala 80:57]
  wire [2:0] _atomics_T_9_opcode = 5'h8 == s2_req_cmd ? 3'h2 : _atomics_T_7_opcode; // @[Mux.scala 80:57]
  wire [2:0] _atomics_T_9_param = 5'h8 == s2_req_cmd ? 3'h4 : _atomics_T_7_param; // @[Mux.scala 80:57]
  wire [3:0] _atomics_T_9_size = 5'h8 == s2_req_cmd ? atomics_a_size : _atomics_T_7_size; // @[Mux.scala 80:57]
  wire  _atomics_T_9_source = 5'h8 == s2_req_cmd ? a_source : _atomics_T_7_source; // @[Mux.scala 80:57]
  wire [31:0] _atomics_T_9_address = 5'h8 == s2_req_cmd ? atomics_a_address : _atomics_T_7_address; // @[Mux.scala 80:57]
  wire [7:0] _atomics_T_9_mask = 5'h8 == s2_req_cmd ? get_mask : _atomics_T_7_mask; // @[Mux.scala 80:57]
  wire [63:0] _atomics_T_9_data = 5'h8 == s2_req_cmd ? pstore1_data : _atomics_T_7_data; // @[Mux.scala 80:57]
  wire [2:0] _atomics_T_11_opcode = 5'hc == s2_req_cmd ? 3'h2 : _atomics_T_9_opcode; // @[Mux.scala 80:57]
  wire [2:0] _atomics_T_11_param = 5'hc == s2_req_cmd ? 3'h0 : _atomics_T_9_param; // @[Mux.scala 80:57]
  wire [3:0] _atomics_T_11_size = 5'hc == s2_req_cmd ? atomics_a_size : _atomics_T_9_size; // @[Mux.scala 80:57]
  wire  _atomics_T_11_source = 5'hc == s2_req_cmd ? a_source : _atomics_T_9_source; // @[Mux.scala 80:57]
  wire [31:0] _atomics_T_11_address = 5'hc == s2_req_cmd ? atomics_a_address : _atomics_T_9_address; // @[Mux.scala 80:57]
  wire [7:0] _atomics_T_11_mask = 5'hc == s2_req_cmd ? get_mask : _atomics_T_9_mask; // @[Mux.scala 80:57]
  wire [63:0] _atomics_T_11_data = 5'hc == s2_req_cmd ? pstore1_data : _atomics_T_9_data; // @[Mux.scala 80:57]
  wire [2:0] _atomics_T_13_opcode = 5'hd == s2_req_cmd ? 3'h2 : _atomics_T_11_opcode; // @[Mux.scala 80:57]
  wire [2:0] _atomics_T_13_param = 5'hd == s2_req_cmd ? 3'h1 : _atomics_T_11_param; // @[Mux.scala 80:57]
  wire [3:0] _atomics_T_13_size = 5'hd == s2_req_cmd ? atomics_a_size : _atomics_T_11_size; // @[Mux.scala 80:57]
  wire  _atomics_T_13_source = 5'hd == s2_req_cmd ? a_source : _atomics_T_11_source; // @[Mux.scala 80:57]
  wire [31:0] _atomics_T_13_address = 5'hd == s2_req_cmd ? atomics_a_address : _atomics_T_11_address; // @[Mux.scala 80:57]
  wire [7:0] _atomics_T_13_mask = 5'hd == s2_req_cmd ? get_mask : _atomics_T_11_mask; // @[Mux.scala 80:57]
  wire [63:0] _atomics_T_13_data = 5'hd == s2_req_cmd ? pstore1_data : _atomics_T_11_data; // @[Mux.scala 80:57]
  wire [2:0] _atomics_T_15_opcode = 5'he == s2_req_cmd ? 3'h2 : _atomics_T_13_opcode; // @[Mux.scala 80:57]
  wire [2:0] _atomics_T_15_param = 5'he == s2_req_cmd ? 3'h2 : _atomics_T_13_param; // @[Mux.scala 80:57]
  wire [3:0] _atomics_T_15_size = 5'he == s2_req_cmd ? atomics_a_size : _atomics_T_13_size; // @[Mux.scala 80:57]
  wire  _atomics_T_15_source = 5'he == s2_req_cmd ? a_source : _atomics_T_13_source; // @[Mux.scala 80:57]
  wire [31:0] _atomics_T_15_address = 5'he == s2_req_cmd ? atomics_a_address : _atomics_T_13_address; // @[Mux.scala 80:57]
  wire [7:0] _atomics_T_15_mask = 5'he == s2_req_cmd ? get_mask : _atomics_T_13_mask; // @[Mux.scala 80:57]
  wire [63:0] _atomics_T_15_data = 5'he == s2_req_cmd ? pstore1_data : _atomics_T_13_data; // @[Mux.scala 80:57]
  wire [2:0] atomics_opcode = 5'hf == s2_req_cmd ? 3'h2 : _atomics_T_15_opcode; // @[Mux.scala 80:57]
  wire [2:0] atomics_param = 5'hf == s2_req_cmd ? 3'h3 : _atomics_T_15_param; // @[Mux.scala 80:57]
  wire [3:0] atomics_size = 5'hf == s2_req_cmd ? atomics_a_size : _atomics_T_15_size; // @[Mux.scala 80:57]
  wire  atomics_source = 5'hf == s2_req_cmd ? a_source : _atomics_T_15_source; // @[Mux.scala 80:57]
  wire [31:0] atomics_address = 5'hf == s2_req_cmd ? atomics_a_address : _atomics_T_15_address; // @[Mux.scala 80:57]
  wire [7:0] atomics_mask = 5'hf == s2_req_cmd ? get_mask : _atomics_T_15_mask; // @[Mux.scala 80:57]
  wire [63:0] atomics_data = 5'hf == s2_req_cmd ? pstore1_data : _atomics_T_15_data; // @[Mux.scala 80:57]
  wire  _tl_out_a_valid_T_6 = (s2_valid_cached_miss & (~release_ack_wait)) & (~s2_victim_dirty); // @[DCache.scala 551:48]
  wire  tl_out_a_valid = s2_valid_uncached_pending | _tl_out_a_valid_T_6; // @[DCache.scala 550:67]
  wire  _tl_out_a_bits_T_3 = ~s2_write; // @[DCache.scala 553:9]
  wire  _tl_out_a_bits_T_5 = ~s2_read; // @[DCache.scala 555:9]
  wire [2:0] _tl_out_a_bits_T_6_opcode = _tl_out_a_bits_T_5 ? 3'h0 : atomics_opcode; // @[DCache.scala 555:8]
  wire [2:0] _tl_out_a_bits_T_6_param = _tl_out_a_bits_T_5 ? 3'h0 : atomics_param; // @[DCache.scala 555:8]
  wire [3:0] _tl_out_a_bits_T_6_size = _tl_out_a_bits_T_5 ? atomics_a_size : atomics_size; // @[DCache.scala 555:8]
  wire  _tl_out_a_bits_T_6_source = ~s2_read ? a_source : atomics_source; // @[DCache.scala 555:8]
  wire [31:0] _tl_out_a_bits_T_6_address = _tl_out_a_bits_T_5 ? atomics_a_address : atomics_address; // @[DCache.scala 555:8]
  wire [7:0] _tl_out_a_bits_T_6_mask = _tl_out_a_bits_T_5 ? get_mask : atomics_mask; // @[DCache.scala 555:8]
  wire [63:0] _tl_out_a_bits_T_6_data = _tl_out_a_bits_T_5 ? pstore1_data : atomics_data; // @[DCache.scala 555:8]
  wire [2:0] _tl_out_a_bits_T_7_opcode = _s2_write_T_1 ? 3'h1 : _tl_out_a_bits_T_6_opcode; // @[DCache.scala 554:8]
  wire [2:0] _tl_out_a_bits_T_7_param = _s2_write_T_1 ? 3'h0 : _tl_out_a_bits_T_6_param; // @[DCache.scala 554:8]
  wire [3:0] _tl_out_a_bits_T_7_size = _s2_write_T_1 ? atomics_a_size : _tl_out_a_bits_T_6_size; // @[DCache.scala 554:8]
  wire  _tl_out_a_bits_T_7_source = _s2_write_T_1 ? a_source : _tl_out_a_bits_T_6_source; // @[DCache.scala 554:8]
  wire [31:0] _tl_out_a_bits_T_7_address = _s2_write_T_1 ? atomics_a_address : _tl_out_a_bits_T_6_address; // @[DCache.scala 554:8]
  wire [7:0] putpartial_mask = a_mask[7:0]; // @[Edges.scala 485:17 Edges.scala 491:15]
  wire [7:0] _tl_out_a_bits_T_7_mask = _s2_write_T_1 ? putpartial_mask : _tl_out_a_bits_T_6_mask; // @[DCache.scala 554:8]
  wire [63:0] _tl_out_a_bits_T_7_data = _s2_write_T_1 ? pstore1_data : _tl_out_a_bits_T_6_data; // @[DCache.scala 554:8]
  wire [2:0] _tl_out_a_bits_T_8_opcode = _tl_out_a_bits_T_3 ? 3'h4 : _tl_out_a_bits_T_7_opcode; // @[DCache.scala 553:8]
  wire [2:0] _tl_out_a_bits_T_8_param = _tl_out_a_bits_T_3 ? 3'h0 : _tl_out_a_bits_T_7_param; // @[DCache.scala 553:8]
  wire [3:0] _tl_out_a_bits_T_8_size = _tl_out_a_bits_T_3 ? atomics_a_size : _tl_out_a_bits_T_7_size; // @[DCache.scala 553:8]
  wire  _tl_out_a_bits_T_8_source = ~s2_write ? a_source : _tl_out_a_bits_T_7_source; // @[DCache.scala 553:8]
  wire [31:0] _tl_out_a_bits_T_8_address = _tl_out_a_bits_T_3 ? atomics_a_address : _tl_out_a_bits_T_7_address; // @[DCache.scala 553:8]
  wire [7:0] _tl_out_a_bits_T_8_mask = _tl_out_a_bits_T_3 ? get_mask : _tl_out_a_bits_T_7_mask; // @[DCache.scala 553:8]
  wire [63:0] _tl_out_a_bits_T_8_data = _tl_out_a_bits_T_3 ? 64'h0 : _tl_out_a_bits_T_7_data; // @[DCache.scala 553:8]
  wire [2:0] tl_out_a_bits_a_param = {{1'd0}, s2_grow_param}; // @[Edges.scala 347:17 Edges.scala 349:15]
  wire [31:0] tl_out_a_bits_a_address = acquire_address[31:0]; // @[Edges.scala 347:17 Edges.scala 352:15]
  wire [1:0] _a_sel_T = 2'h1 << a_source; // @[OneHot.scala 65:12]
  wire  a_sel = _a_sel_T[1]; // @[DCache.scala 574:66]
  wire  _T_228 = auto_out_a_ready & tl_out_a_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_143 = a_sel | uncachedInFlight_0; // @[DCache.scala 578:18 DCache.scala 579:13 DCache.scala 206:33]
  wire  _GEN_155 = s2_uncached ? _GEN_143 : uncachedInFlight_0; // @[DCache.scala 576:24 DCache.scala 206:33]
  wire  _GEN_167 = s2_uncached ? cached_grant_wait : 1'h1; // @[DCache.scala 576:24 DCache.scala 196:30 DCache.scala 585:25]
  wire  _GEN_168 = _T_228 ? _GEN_155 : uncachedInFlight_0; // @[DCache.scala 575:26 DCache.scala 206:33]
  wire  _GEN_180 = _T_228 ? _GEN_167 : cached_grant_wait; // @[DCache.scala 575:26 DCache.scala 196:30]
  wire [26:0] _beats1_decode_T_1 = 27'hfff << auto_out_d_bits_size; // @[package.scala 212:77]
  wire [11:0] _beats1_decode_T_3 = ~(_beats1_decode_T_1[11:0]); // @[package.scala 212:46]
  wire [8:0] beats1_decode = _beats1_decode_T_3[11:3]; // @[Edges.scala 221:59]
  wire  beats1_opdata = auto_out_d_bits_opcode[0]; // @[Edges.scala 107:36]
  wire [8:0] beats1 = beats1_opdata ? beats1_decode : 9'h0; // @[Edges.scala 222:14]
  wire [8:0] counter1 = counter - 9'h1; // @[Edges.scala 231:28]
  wire  d_last = (counter == 9'h1) | (beats1 == 9'h0); // @[Edges.scala 233:37]
  wire  d_done = d_last & _T_236; // @[Edges.scala 234:22]
  wire [8:0] _count_T = ~counter1; // @[Edges.scala 235:27]
  wire [8:0] count = beats1 & _count_T; // @[Edges.scala 235:25]
  wire [11:0] d_address_inc = {count, 3'h0}; // @[Edges.scala 270:29]
  wire  _tl_d_data_encoded_T_4 = ~grantIsUncached; // @[DCache.scala 606:129]
  wire  grantIsVoluntary = auto_out_d_bits_opcode == 3'h6; // @[DCache.scala 608:32]
  wire [2:0] _blockProbeAfterGrantCount_T_1 = blockProbeAfterGrantCount - 3'h1; // @[DCache.scala 612:97]
  wire [2:0] _GEN_182 = _block_probe_for_core_progress_T ? _blockProbeAfterGrantCount_T_1 : blockProbeAfterGrantCount; // @[DCache.scala 612:40 DCache.scala 612:68 DCache.scala 611:38]
  wire [1:0] _uncachedRespIdxOH_T = 2'h1 << auto_out_d_bits_source; // @[OneHot.scala 65:12]
  wire  uncachedRespIdxOH = _uncachedRespIdxOH_T[1]; // @[DCache.scala 615:90]
  wire  _T_241 = uncachedRespIdxOH & d_last; // @[DCache.scala 629:17]
  wire  _GEN_187 = _T_241 ? 1'h0 : _GEN_168; // @[DCache.scala 629:28 DCache.scala 631:13]
  wire [31:0] dontCareBits = {s1_paddr[31:3], 3'h0}; // @[DCache.scala 644:55]
  wire [31:0] _GEN_392 = {{29'd0}, uncachedReqs_0_addr[2:0]}; // @[DCache.scala 645:26]
  wire [31:0] _s2_req_addr_T_1 = dontCareBits | _GEN_392; // @[DCache.scala 645:26]
  wire  _GEN_195 = grantIsVoluntary ? 1'h0 : release_ack_wait; // @[DCache.scala 650:36 DCache.scala 652:24 DCache.scala 197:29]
  wire  _GEN_204 = grantIsUncached ? release_ack_wait : _GEN_195; // @[DCache.scala 627:35 DCache.scala 197:29]
  wire  _GEN_208 = grantIsCached & d_last; // @[DCache.scala 618:26 Replacement.scala 37:11]
  wire  _GEN_217 = grantIsCached ? release_ack_wait : _GEN_204; // @[DCache.scala 618:26 DCache.scala 197:29]
  wire  _GEN_230 = _T_236 ? _GEN_217 : release_ack_wait; // @[DCache.scala 617:26 DCache.scala 197:29]
  wire  _tl_out_e_valid_T_2 = ((auto_out_d_valid & d_first) & grantIsCached) & canAcceptCachedGrant; // @[DCache.scala 657:64]
  wire  tl_out__e_valid = _T_257 ? 1'h0 : _tl_out_e_valid_T_2; // @[DCache.scala 665:51 DCache.scala 666:20 DCache.scala 657:18]
  wire  _T_248 = auto_out_e_ready & tl_out__e_valid; // @[Decoupled.scala 40:37]
  wire  _dataArb_io_in_1_valid_T_1 = (auto_out_d_valid & grantIsRefill) & canAcceptCachedGrant; // @[DCache.scala 664:61]
  wire [39:0] _dataArb_io_in_1_bits_addr_T_1 = {s2_vaddr[39:6], 6'h0}; // @[DCache.scala 671:57]
  wire [39:0] _GEN_393 = {{28'd0}, d_address_inc}; // @[DCache.scala 671:67]
  wire [39:0] _dataArb_io_in_1_bits_addr_T_2 = _dataArb_io_in_1_bits_addr_T_1 | _GEN_393; // @[DCache.scala 671:67]
  wire [3:0] _metaArb_io_in_3_bits_data_T_1 = {s2_write,c_cat_left,auto_out_d_bits_param}; // @[Cat.scala 29:58]
  wire [1:0] _metaArb_io_in_3_bits_data_T_7 = 4'h1 == _metaArb_io_in_3_bits_data_T_1 ? 2'h1 : 2'h0; // @[Mux.scala 80:57]
  wire [1:0] _metaArb_io_in_3_bits_data_T_9 = 4'h0 == _metaArb_io_in_3_bits_data_T_1 ? 2'h2 :
    _metaArb_io_in_3_bits_data_T_7; // @[Mux.scala 80:57]
  wire [1:0] _metaArb_io_in_3_bits_data_T_11 = 4'h4 == _metaArb_io_in_3_bits_data_T_1 ? 2'h2 :
    _metaArb_io_in_3_bits_data_T_9; // @[Mux.scala 80:57]
  wire [1:0] metaArb_io_in_3_bits_data_meta_state = 4'hc == _metaArb_io_in_3_bits_data_T_1 ? 2'h3 :
    _metaArb_io_in_3_bits_data_T_11; // @[Mux.scala 80:57]
  wire  _GEN_233 = auto_out_d_valid ? 1'h0 : _GEN_31; // @[DCache.scala 698:29 DCache.scala 699:26]
  wire  _GEN_234 = auto_out_d_valid | _dataArb_io_in_1_valid_T_1; // @[DCache.scala 698:29 DCache.scala 700:32 DCache.scala 664:26]
  wire  _GEN_235 = auto_out_d_valid ? 1'h0 : 1'h1; // @[DCache.scala 698:29 DCache.scala 701:37 DCache.scala 670:33]
  wire  _metaArb_io_in_6_valid_T_2 = auto_out_b_valid & ((~block_probe_for_core_progress) | lrscBackingOff); // @[DCache.scala 712:44]
  wire [7:0] metaArb_io_in_6_bits_addr_right = io_cpu_req_bits_addr[39:32]; // @[DCache.scala 716:58]
  wire [39:0] _metaArb_io_in_6_bits_addr_T = {metaArb_io_in_6_bits_addr_right,auto_out_b_bits_address}; // @[Cat.scala 29:58]
  wire [8:0] counter1_1 = counter_1 - 9'h1; // @[Edges.scala 231:28]
  wire [8:0] _count_T_1 = ~counter1_1; // @[Edges.scala 235:27]
  wire [8:0] c_count = beats1_1 & _count_T_1; // @[Edges.scala 235:25]
  reg  s1_release_data_valid; // @[DCache.scala 723:34]
  wire  releaseRejected = s2_release_data_valid & (~_T_262); // @[DCache.scala 725:44]
  wire [9:0] _releaseDataBeat_T = {1'h0,c_count}; // @[Cat.scala 29:58]
  wire [1:0] _releaseDataBeat_T_1 = {1'h0,s2_release_data_valid}; // @[Cat.scala 29:58]
  wire [1:0] _GEN_394 = {{1'd0}, s1_release_data_valid}; // @[DCache.scala 726:101]
  wire [1:0] _releaseDataBeat_T_3 = _GEN_394 + _releaseDataBeat_T_1; // @[DCache.scala 726:101]
  wire [1:0] _releaseDataBeat_T_4 = releaseRejected ? 2'h0 : _releaseDataBeat_T_3; // @[DCache.scala 726:52]
  wire [9:0] _GEN_395 = {{8'd0}, _releaseDataBeat_T_4}; // @[DCache.scala 726:47]
  wire [9:0] releaseDataBeat = _releaseDataBeat_T + _GEN_395; // @[DCache.scala 726:47]
  wire  discard_line = s2_valid_flush_line & (s2_req_size[1]); // @[DCache.scala 740:46]
  wire  _release_state_T_1 = s2_victim_dirty & (~discard_line); // @[DCache.scala 741:44]
  wire [2:0] _release_state_T_2 = _release_state_T_1 ? 3'h1 : 3'h6; // @[DCache.scala 741:27]
  wire [5:0] probe_bits_left = s2_req_addr[11:6]; // @[DCache.scala 742:76]
  wire [25:0] _probe_bits_T_1 = {s2_victim_tag,probe_bits_left}; // @[Cat.scala 29:58]
  wire [31:0] res_2_address = {_probe_bits_T_1, 6'h0}; // @[DCache.scala 742:96]
  wire [2:0] _GEN_243 = s2_want_victimize ? _release_state_T_2 : release_state; // @[DCache.scala 738:25 DCache.scala 741:21 DCache.scala 199:26]
  wire [2:0] _release_state_T_3 = releaseDone ? 3'h7 : 3'h3; // @[DCache.scala 753:29]
  wire [2:0] _release_state_T_4 = releaseDone ? 3'h0 : 3'h5; // @[DCache.scala 757:29]
  wire [2:0] _GEN_254 = _T_268 ? s2_report_param : 3'h5; // @[DCache.scala 750:45 DCache.scala 752:23 DCache.scala 733:17]
  wire [2:0] _GEN_260 = _T_268 ? _release_state_T_3 : _release_state_T_4; // @[DCache.scala 750:45 DCache.scala 753:23 DCache.scala 757:23]
  wire [2:0] _GEN_262 = s2_prb_ack_data ? 3'h2 : _GEN_260; // @[DCache.scala 748:36 DCache.scala 749:23]
  wire [2:0] _GEN_265 = s2_prb_ack_data ? 3'h5 : _GEN_254; // @[DCache.scala 748:36 DCache.scala 733:17]
  wire [2:0] _GEN_283 = s2_probe ? _GEN_262 : _GEN_243; // @[DCache.scala 744:21]
  wire [2:0] _GEN_286 = s2_probe ? _GEN_265 : 3'h5; // @[DCache.scala 744:21 DCache.scala 733:17]
  wire  _T_269 = release_state == 3'h4; // @[DCache.scala 761:25]
  wire [39:0] _metaArb_io_in_6_bits_addr_T_1 = {metaArb_io_in_6_bits_addr_right,probe_bits_address}; // @[Cat.scala 29:58]
  wire [2:0] _GEN_293 = metaArb_io_in_6_ready ? 3'h0 : _GEN_283; // @[DCache.scala 765:37 DCache.scala 766:23]
  wire  _GEN_294 = metaArb_io_in_6_ready | s1_probe_x12; // @[DCache.scala 765:37 DCache.scala 767:18 DCache.scala 160:21]
  wire [2:0] _GEN_298 = _T_269 ? _GEN_293 : _GEN_283; // @[DCache.scala 761:44]
  wire [2:0] _GEN_300 = releaseDone ? 3'h0 : _GEN_298; // @[DCache.scala 772:26 DCache.scala 772:42]
  wire [2:0] _GEN_302 = _T_270 ? _GEN_300 : _GEN_298; // @[DCache.scala 770:47]
  wire [2:0] _GEN_303 = releaseDone ? 3'h7 : _GEN_302; // @[DCache.scala 777:26 DCache.scala 777:42]
  wire [2:0] _GEN_306 = _T_271 ? s2_report_param : _GEN_286; // @[DCache.scala 774:48 DCache.scala 776:21]
  wire [2:0] _GEN_312 = _T_271 ? _GEN_303 : _GEN_302; // @[DCache.scala 774:48]
  wire [2:0] _GEN_313 = releaseDone ? 3'h7 : _GEN_312; // @[DCache.scala 781:26 DCache.scala 781:42]
  wire [2:0] _GEN_315 = _T_272 ? s2_report_param : _GEN_306; // @[DCache.scala 779:48 DCache.scala 780:21]
  wire [2:0] _GEN_321 = _T_272 ? _GEN_313 : _GEN_312; // @[DCache.scala 779:48]
  wire  _T_277 = _T_262 & c_first; // @[DCache.scala 792:29]
  wire  _GEN_323 = _T_277 | _GEN_230; // @[DCache.scala 792:41 DCache.scala 793:26]
  wire [1:0] newCoh_state = _T_275 ? voluntaryNewCoh_state : probeNewCoh_state; // @[DCache.scala 783:81 DCache.scala 789:14]
  wire [11:0] _dataArb_io_in_2_bits_addr_T_1 = {probe_bits_address[11:6], 6'h0}; // @[DCache.scala 806:55]
  wire [5:0] _dataArb_io_in_2_bits_addr_T_3 = {releaseDataBeat[2:0], 3'h0}; // @[DCache.scala 806:117]
  wire [11:0] _GEN_397 = {{6'd0}, _dataArb_io_in_2_bits_addr_T_3}; // @[DCache.scala 806:72]
  wire  _metaArb_io_in_4_valid_T_1 = release_state == 3'h7; // @[package.scala 15:47]
  wire [11:0] metaArb_io_in_4_bits_addr_left = probe_bits_address[11:0]; // @[DCache.scala 814:90]
  wire [19:0] metaArb_io_in_4_bits_data_meta_tag = probe_bits_address[31:12]; // @[DCache.scala 815:78]
  wire  _T_278 = metaArb_io_in_4_ready & metaArb_io_in_4_valid; // @[Decoupled.scala 40:37]
  reg  io_cpu_s2_xcpt_REG; // @[DCache.scala 832:32]
  reg  doUncachedResp; // @[DCache.scala 847:27]
  wire [31:0] io_cpu_resp_bits_data_shifted = get_get_mask_bit ? s2_data_corrected[63:32] : s2_data_corrected[31:0]; // @[AMOALU.scala 39:24]
  wire  _io_cpu_resp_bits_data_T_3 = s2_req_signed & (io_cpu_resp_bits_data_shifted[31]); // @[AMOALU.scala 42:76]
  wire [31:0] _io_cpu_resp_bits_data_T_5 = _io_cpu_resp_bits_data_T_3 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] io_cpu_resp_bits_data_right = s2_req_size == 2'h2 ? _io_cpu_resp_bits_data_T_5 : s2_data_corrected[63:32]; // @[AMOALU.scala 42:20]
  wire [63:0] _io_cpu_resp_bits_data_T_7 = {io_cpu_resp_bits_data_right,io_cpu_resp_bits_data_shifted}; // @[Cat.scala 29:58]
  wire [15:0] io_cpu_resp_bits_data_shifted_1 = get_get_mask_bit_1 ? _io_cpu_resp_bits_data_T_7[31:16] :
    _io_cpu_resp_bits_data_T_7[15:0]; // @[AMOALU.scala 39:24]
  wire  _io_cpu_resp_bits_data_T_11 = s2_req_signed & (io_cpu_resp_bits_data_shifted_1[15]); // @[AMOALU.scala 42:76]
  wire [47:0] _io_cpu_resp_bits_data_T_13 = _io_cpu_resp_bits_data_T_11 ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 72:12]
  wire [47:0] io_cpu_resp_bits_data_right_1 = s2_req_size == 2'h1 ? _io_cpu_resp_bits_data_T_13 :
    _io_cpu_resp_bits_data_T_7[63:16]; // @[AMOALU.scala 42:20]
  wire [63:0] _io_cpu_resp_bits_data_T_15 = {io_cpu_resp_bits_data_right_1,io_cpu_resp_bits_data_shifted_1}; // @[Cat.scala 29:58]
  wire [7:0] io_cpu_resp_bits_data_shifted_2 = get_get_mask_bit_2 ? _io_cpu_resp_bits_data_T_15[15:8] :
    _io_cpu_resp_bits_data_T_15[7:0]; // @[AMOALU.scala 39:24]
  wire [7:0] io_cpu_resp_bits_data_left_2 = _s2_write_T_3 ? 8'h0 : io_cpu_resp_bits_data_shifted_2; // @[AMOALU.scala 41:23]
  wire  _io_cpu_resp_bits_data_T_17 = (s2_req_size == 2'h0) | _s2_write_T_3; // @[AMOALU.scala 42:38]
  wire  _io_cpu_resp_bits_data_T_19 = s2_req_signed & (io_cpu_resp_bits_data_left_2[7]); // @[AMOALU.scala 42:76]
  wire [55:0] _io_cpu_resp_bits_data_T_21 = _io_cpu_resp_bits_data_T_19 ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 72:12]
  wire [55:0] io_cpu_resp_bits_data_right_2 = _io_cpu_resp_bits_data_T_17 ? _io_cpu_resp_bits_data_T_21 :
    _io_cpu_resp_bits_data_T_15[63:8]; // @[AMOALU.scala 42:20]
  wire [63:0] _io_cpu_resp_bits_data_T_23 = {io_cpu_resp_bits_data_right_2,io_cpu_resp_bits_data_left_2}; // @[Cat.scala 29:58]
  wire [63:0] _GEN_398 = {{63'd0}, s2_sc_fail}; // @[DCache.scala 873:41]
  reg  resetting; // @[DCache.scala 906:26]
  reg  REG; // @[DCache.scala 908:18]
  wire  _GEN_341 = REG | resetting; // @[DCache.scala 908:27 DCache.scala 908:39 DCache.scala 906:26]
  reg [7:0] flushCounter; // @[DCache.scala 909:25]
  wire [8:0] flushCounterNext = flushCounter + 8'h1; // @[DCache.scala 910:39]
  wire  flushDone = (flushCounterNext[8:6]) == 3'h4; // @[DCache.scala 911:57]
  wire [11:0] metaArb_io_in_5_bits_addr_left = {metaArb_io_in_5_bits_idx, 6'h0}; // @[DCache.scala 919:98]
  wire [8:0] _GEN_343 = resetting ? flushCounterNext : {{1'd0}, flushCounter}; // @[DCache.scala 952:20 DCache.scala 953:18 DCache.scala 909:25]
  reg [8:0] io_cpu_perf_release_counter; // @[Edges.scala 230:27]
  wire [8:0] io_cpu_perf_release_counter1 = io_cpu_perf_release_counter - 9'h1; // @[Edges.scala 231:28]
  wire  io_cpu_perf_release_first = io_cpu_perf_release_counter == 9'h0; // @[Edges.scala 232:25]
  wire  io_cpu_perf_release_last = (io_cpu_perf_release_counter == 9'h1) | (beats1_1 == 9'h0); // @[Edges.scala 233:37]
  wire  _T_294 = ~grantIsCached; // @[DCache.scala 1028:35]
  wire  _GEN_404 = _T_236 & _T_294; // @[DCache.scala 630:17]
  OptimizationBarrier tlb_mpu_ppn_data_barrier ( // @[package.scala 236:25]
    .io_x_ppn(tlb_mpu_ppn_data_barrier_io_x_ppn),
    .io_x_u(tlb_mpu_ppn_data_barrier_io_x_u),
    .io_x_ae(tlb_mpu_ppn_data_barrier_io_x_ae),
    .io_x_sw(tlb_mpu_ppn_data_barrier_io_x_sw),
    .io_x_sx(tlb_mpu_ppn_data_barrier_io_x_sx),
    .io_x_sr(tlb_mpu_ppn_data_barrier_io_x_sr),
    .io_x_pw(tlb_mpu_ppn_data_barrier_io_x_pw),
    .io_x_px(tlb_mpu_ppn_data_barrier_io_x_px),
    .io_x_pr(tlb_mpu_ppn_data_barrier_io_x_pr),
    .io_x_ppp(tlb_mpu_ppn_data_barrier_io_x_ppp),
    .io_x_pal(tlb_mpu_ppn_data_barrier_io_x_pal),
    .io_x_paa(tlb_mpu_ppn_data_barrier_io_x_paa),
    .io_x_eff(tlb_mpu_ppn_data_barrier_io_x_eff),
    .io_x_c(tlb_mpu_ppn_data_barrier_io_x_c),
    .io_y_ppn(tlb_mpu_ppn_data_barrier_io_y_ppn),
    .io_y_u(tlb_mpu_ppn_data_barrier_io_y_u),
    .io_y_ae(tlb_mpu_ppn_data_barrier_io_y_ae),
    .io_y_sw(tlb_mpu_ppn_data_barrier_io_y_sw),
    .io_y_sx(tlb_mpu_ppn_data_barrier_io_y_sx),
    .io_y_sr(tlb_mpu_ppn_data_barrier_io_y_sr),
    .io_y_pw(tlb_mpu_ppn_data_barrier_io_y_pw),
    .io_y_px(tlb_mpu_ppn_data_barrier_io_y_px),
    .io_y_pr(tlb_mpu_ppn_data_barrier_io_y_pr),
    .io_y_ppp(tlb_mpu_ppn_data_barrier_io_y_ppp),
    .io_y_pal(tlb_mpu_ppn_data_barrier_io_y_pal),
    .io_y_paa(tlb_mpu_ppn_data_barrier_io_y_paa),
    .io_y_eff(tlb_mpu_ppn_data_barrier_io_y_eff),
    .io_y_c(tlb_mpu_ppn_data_barrier_io_y_c)
  );
  PMPChecker tlb_pmp ( // @[TLB.scala 190:19]
    .io_prv(tlb_pmp_io_prv),
    .io_pmp_0_cfg_l(tlb_pmp_io_pmp_0_cfg_l),
    .io_pmp_0_cfg_a(tlb_pmp_io_pmp_0_cfg_a),
    .io_pmp_0_cfg_x(tlb_pmp_io_pmp_0_cfg_x),
    .io_pmp_0_cfg_w(tlb_pmp_io_pmp_0_cfg_w),
    .io_pmp_0_cfg_r(tlb_pmp_io_pmp_0_cfg_r),
    .io_pmp_0_addr(tlb_pmp_io_pmp_0_addr),
    .io_pmp_0_mask(tlb_pmp_io_pmp_0_mask),
    .io_pmp_1_cfg_l(tlb_pmp_io_pmp_1_cfg_l),
    .io_pmp_1_cfg_a(tlb_pmp_io_pmp_1_cfg_a),
    .io_pmp_1_cfg_x(tlb_pmp_io_pmp_1_cfg_x),
    .io_pmp_1_cfg_w(tlb_pmp_io_pmp_1_cfg_w),
    .io_pmp_1_cfg_r(tlb_pmp_io_pmp_1_cfg_r),
    .io_pmp_1_addr(tlb_pmp_io_pmp_1_addr),
    .io_pmp_1_mask(tlb_pmp_io_pmp_1_mask),
    .io_pmp_2_cfg_l(tlb_pmp_io_pmp_2_cfg_l),
    .io_pmp_2_cfg_a(tlb_pmp_io_pmp_2_cfg_a),
    .io_pmp_2_cfg_x(tlb_pmp_io_pmp_2_cfg_x),
    .io_pmp_2_cfg_w(tlb_pmp_io_pmp_2_cfg_w),
    .io_pmp_2_cfg_r(tlb_pmp_io_pmp_2_cfg_r),
    .io_pmp_2_addr(tlb_pmp_io_pmp_2_addr),
    .io_pmp_2_mask(tlb_pmp_io_pmp_2_mask),
    .io_pmp_3_cfg_l(tlb_pmp_io_pmp_3_cfg_l),
    .io_pmp_3_cfg_a(tlb_pmp_io_pmp_3_cfg_a),
    .io_pmp_3_cfg_x(tlb_pmp_io_pmp_3_cfg_x),
    .io_pmp_3_cfg_w(tlb_pmp_io_pmp_3_cfg_w),
    .io_pmp_3_cfg_r(tlb_pmp_io_pmp_3_cfg_r),
    .io_pmp_3_addr(tlb_pmp_io_pmp_3_addr),
    .io_pmp_3_mask(tlb_pmp_io_pmp_3_mask),
    .io_pmp_4_cfg_l(tlb_pmp_io_pmp_4_cfg_l),
    .io_pmp_4_cfg_a(tlb_pmp_io_pmp_4_cfg_a),
    .io_pmp_4_cfg_x(tlb_pmp_io_pmp_4_cfg_x),
    .io_pmp_4_cfg_w(tlb_pmp_io_pmp_4_cfg_w),
    .io_pmp_4_cfg_r(tlb_pmp_io_pmp_4_cfg_r),
    .io_pmp_4_addr(tlb_pmp_io_pmp_4_addr),
    .io_pmp_4_mask(tlb_pmp_io_pmp_4_mask),
    .io_pmp_5_cfg_l(tlb_pmp_io_pmp_5_cfg_l),
    .io_pmp_5_cfg_a(tlb_pmp_io_pmp_5_cfg_a),
    .io_pmp_5_cfg_x(tlb_pmp_io_pmp_5_cfg_x),
    .io_pmp_5_cfg_w(tlb_pmp_io_pmp_5_cfg_w),
    .io_pmp_5_cfg_r(tlb_pmp_io_pmp_5_cfg_r),
    .io_pmp_5_addr(tlb_pmp_io_pmp_5_addr),
    .io_pmp_5_mask(tlb_pmp_io_pmp_5_mask),
    .io_pmp_6_cfg_l(tlb_pmp_io_pmp_6_cfg_l),
    .io_pmp_6_cfg_a(tlb_pmp_io_pmp_6_cfg_a),
    .io_pmp_6_cfg_x(tlb_pmp_io_pmp_6_cfg_x),
    .io_pmp_6_cfg_w(tlb_pmp_io_pmp_6_cfg_w),
    .io_pmp_6_cfg_r(tlb_pmp_io_pmp_6_cfg_r),
    .io_pmp_6_addr(tlb_pmp_io_pmp_6_addr),
    .io_pmp_6_mask(tlb_pmp_io_pmp_6_mask),
    .io_pmp_7_cfg_l(tlb_pmp_io_pmp_7_cfg_l),
    .io_pmp_7_cfg_a(tlb_pmp_io_pmp_7_cfg_a),
    .io_pmp_7_cfg_x(tlb_pmp_io_pmp_7_cfg_x),
    .io_pmp_7_cfg_w(tlb_pmp_io_pmp_7_cfg_w),
    .io_pmp_7_cfg_r(tlb_pmp_io_pmp_7_cfg_r),
    .io_pmp_7_addr(tlb_pmp_io_pmp_7_addr),
    .io_pmp_7_mask(tlb_pmp_io_pmp_7_mask),
    .io_addr(tlb_pmp_io_addr),
    .io_size(tlb_pmp_io_size),
    .io_r(tlb_pmp_io_r),
    .io_w(tlb_pmp_io_w),
    .io_x(tlb_pmp_io_x)
  );
  OptimizationBarrier tlb_ppn_data_barrier ( // @[package.scala 236:25]
    .io_x_ppn(tlb_ppn_data_barrier_io_x_ppn),
    .io_x_u(tlb_ppn_data_barrier_io_x_u),
    .io_x_ae(tlb_ppn_data_barrier_io_x_ae),
    .io_x_sw(tlb_ppn_data_barrier_io_x_sw),
    .io_x_sx(tlb_ppn_data_barrier_io_x_sx),
    .io_x_sr(tlb_ppn_data_barrier_io_x_sr),
    .io_x_pw(tlb_ppn_data_barrier_io_x_pw),
    .io_x_px(tlb_ppn_data_barrier_io_x_px),
    .io_x_pr(tlb_ppn_data_barrier_io_x_pr),
    .io_x_ppp(tlb_ppn_data_barrier_io_x_ppp),
    .io_x_pal(tlb_ppn_data_barrier_io_x_pal),
    .io_x_paa(tlb_ppn_data_barrier_io_x_paa),
    .io_x_eff(tlb_ppn_data_barrier_io_x_eff),
    .io_x_c(tlb_ppn_data_barrier_io_x_c),
    .io_y_ppn(tlb_ppn_data_barrier_io_y_ppn),
    .io_y_u(tlb_ppn_data_barrier_io_y_u),
    .io_y_ae(tlb_ppn_data_barrier_io_y_ae),
    .io_y_sw(tlb_ppn_data_barrier_io_y_sw),
    .io_y_sx(tlb_ppn_data_barrier_io_y_sx),
    .io_y_sr(tlb_ppn_data_barrier_io_y_sr),
    .io_y_pw(tlb_ppn_data_barrier_io_y_pw),
    .io_y_px(tlb_ppn_data_barrier_io_y_px),
    .io_y_pr(tlb_ppn_data_barrier_io_y_pr),
    .io_y_ppp(tlb_ppn_data_barrier_io_y_ppp),
    .io_y_pal(tlb_ppn_data_barrier_io_y_pal),
    .io_y_paa(tlb_ppn_data_barrier_io_y_paa),
    .io_y_eff(tlb_ppn_data_barrier_io_y_eff),
    .io_y_c(tlb_ppn_data_barrier_io_y_c)
  );
  OptimizationBarrier tlb_ppn_data_barrier_1 ( // @[package.scala 236:25]
    .io_x_ppn(tlb_ppn_data_barrier_1_io_x_ppn),
    .io_x_u(tlb_ppn_data_barrier_1_io_x_u),
    .io_x_ae(tlb_ppn_data_barrier_1_io_x_ae),
    .io_x_sw(tlb_ppn_data_barrier_1_io_x_sw),
    .io_x_sx(tlb_ppn_data_barrier_1_io_x_sx),
    .io_x_sr(tlb_ppn_data_barrier_1_io_x_sr),
    .io_x_pw(tlb_ppn_data_barrier_1_io_x_pw),
    .io_x_px(tlb_ppn_data_barrier_1_io_x_px),
    .io_x_pr(tlb_ppn_data_barrier_1_io_x_pr),
    .io_x_ppp(tlb_ppn_data_barrier_1_io_x_ppp),
    .io_x_pal(tlb_ppn_data_barrier_1_io_x_pal),
    .io_x_paa(tlb_ppn_data_barrier_1_io_x_paa),
    .io_x_eff(tlb_ppn_data_barrier_1_io_x_eff),
    .io_x_c(tlb_ppn_data_barrier_1_io_x_c),
    .io_y_ppn(tlb_ppn_data_barrier_1_io_y_ppn),
    .io_y_u(tlb_ppn_data_barrier_1_io_y_u),
    .io_y_ae(tlb_ppn_data_barrier_1_io_y_ae),
    .io_y_sw(tlb_ppn_data_barrier_1_io_y_sw),
    .io_y_sx(tlb_ppn_data_barrier_1_io_y_sx),
    .io_y_sr(tlb_ppn_data_barrier_1_io_y_sr),
    .io_y_pw(tlb_ppn_data_barrier_1_io_y_pw),
    .io_y_px(tlb_ppn_data_barrier_1_io_y_px),
    .io_y_pr(tlb_ppn_data_barrier_1_io_y_pr),
    .io_y_ppp(tlb_ppn_data_barrier_1_io_y_ppp),
    .io_y_pal(tlb_ppn_data_barrier_1_io_y_pal),
    .io_y_paa(tlb_ppn_data_barrier_1_io_y_paa),
    .io_y_eff(tlb_ppn_data_barrier_1_io_y_eff),
    .io_y_c(tlb_ppn_data_barrier_1_io_y_c)
  );
  OptimizationBarrier tlb_ppn_data_barrier_2 ( // @[package.scala 236:25]
    .io_x_ppn(tlb_ppn_data_barrier_2_io_x_ppn),
    .io_x_u(tlb_ppn_data_barrier_2_io_x_u),
    .io_x_ae(tlb_ppn_data_barrier_2_io_x_ae),
    .io_x_sw(tlb_ppn_data_barrier_2_io_x_sw),
    .io_x_sx(tlb_ppn_data_barrier_2_io_x_sx),
    .io_x_sr(tlb_ppn_data_barrier_2_io_x_sr),
    .io_x_pw(tlb_ppn_data_barrier_2_io_x_pw),
    .io_x_px(tlb_ppn_data_barrier_2_io_x_px),
    .io_x_pr(tlb_ppn_data_barrier_2_io_x_pr),
    .io_x_ppp(tlb_ppn_data_barrier_2_io_x_ppp),
    .io_x_pal(tlb_ppn_data_barrier_2_io_x_pal),
    .io_x_paa(tlb_ppn_data_barrier_2_io_x_paa),
    .io_x_eff(tlb_ppn_data_barrier_2_io_x_eff),
    .io_x_c(tlb_ppn_data_barrier_2_io_x_c),
    .io_y_ppn(tlb_ppn_data_barrier_2_io_y_ppn),
    .io_y_u(tlb_ppn_data_barrier_2_io_y_u),
    .io_y_ae(tlb_ppn_data_barrier_2_io_y_ae),
    .io_y_sw(tlb_ppn_data_barrier_2_io_y_sw),
    .io_y_sx(tlb_ppn_data_barrier_2_io_y_sx),
    .io_y_sr(tlb_ppn_data_barrier_2_io_y_sr),
    .io_y_pw(tlb_ppn_data_barrier_2_io_y_pw),
    .io_y_px(tlb_ppn_data_barrier_2_io_y_px),
    .io_y_pr(tlb_ppn_data_barrier_2_io_y_pr),
    .io_y_ppp(tlb_ppn_data_barrier_2_io_y_ppp),
    .io_y_pal(tlb_ppn_data_barrier_2_io_y_pal),
    .io_y_paa(tlb_ppn_data_barrier_2_io_y_paa),
    .io_y_eff(tlb_ppn_data_barrier_2_io_y_eff),
    .io_y_c(tlb_ppn_data_barrier_2_io_y_c)
  );
  OptimizationBarrier tlb_ppn_data_barrier_3 ( // @[package.scala 236:25]
    .io_x_ppn(tlb_ppn_data_barrier_3_io_x_ppn),
    .io_x_u(tlb_ppn_data_barrier_3_io_x_u),
    .io_x_ae(tlb_ppn_data_barrier_3_io_x_ae),
    .io_x_sw(tlb_ppn_data_barrier_3_io_x_sw),
    .io_x_sx(tlb_ppn_data_barrier_3_io_x_sx),
    .io_x_sr(tlb_ppn_data_barrier_3_io_x_sr),
    .io_x_pw(tlb_ppn_data_barrier_3_io_x_pw),
    .io_x_px(tlb_ppn_data_barrier_3_io_x_px),
    .io_x_pr(tlb_ppn_data_barrier_3_io_x_pr),
    .io_x_ppp(tlb_ppn_data_barrier_3_io_x_ppp),
    .io_x_pal(tlb_ppn_data_barrier_3_io_x_pal),
    .io_x_paa(tlb_ppn_data_barrier_3_io_x_paa),
    .io_x_eff(tlb_ppn_data_barrier_3_io_x_eff),
    .io_x_c(tlb_ppn_data_barrier_3_io_x_c),
    .io_y_ppn(tlb_ppn_data_barrier_3_io_y_ppn),
    .io_y_u(tlb_ppn_data_barrier_3_io_y_u),
    .io_y_ae(tlb_ppn_data_barrier_3_io_y_ae),
    .io_y_sw(tlb_ppn_data_barrier_3_io_y_sw),
    .io_y_sx(tlb_ppn_data_barrier_3_io_y_sx),
    .io_y_sr(tlb_ppn_data_barrier_3_io_y_sr),
    .io_y_pw(tlb_ppn_data_barrier_3_io_y_pw),
    .io_y_px(tlb_ppn_data_barrier_3_io_y_px),
    .io_y_pr(tlb_ppn_data_barrier_3_io_y_pr),
    .io_y_ppp(tlb_ppn_data_barrier_3_io_y_ppp),
    .io_y_pal(tlb_ppn_data_barrier_3_io_y_pal),
    .io_y_paa(tlb_ppn_data_barrier_3_io_y_paa),
    .io_y_eff(tlb_ppn_data_barrier_3_io_y_eff),
    .io_y_c(tlb_ppn_data_barrier_3_io_y_c)
  );
  OptimizationBarrier tlb_ppn_data_barrier_4 ( // @[package.scala 236:25]
    .io_x_ppn(tlb_ppn_data_barrier_4_io_x_ppn),
    .io_x_u(tlb_ppn_data_barrier_4_io_x_u),
    .io_x_ae(tlb_ppn_data_barrier_4_io_x_ae),
    .io_x_sw(tlb_ppn_data_barrier_4_io_x_sw),
    .io_x_sx(tlb_ppn_data_barrier_4_io_x_sx),
    .io_x_sr(tlb_ppn_data_barrier_4_io_x_sr),
    .io_x_pw(tlb_ppn_data_barrier_4_io_x_pw),
    .io_x_px(tlb_ppn_data_barrier_4_io_x_px),
    .io_x_pr(tlb_ppn_data_barrier_4_io_x_pr),
    .io_x_ppp(tlb_ppn_data_barrier_4_io_x_ppp),
    .io_x_pal(tlb_ppn_data_barrier_4_io_x_pal),
    .io_x_paa(tlb_ppn_data_barrier_4_io_x_paa),
    .io_x_eff(tlb_ppn_data_barrier_4_io_x_eff),
    .io_x_c(tlb_ppn_data_barrier_4_io_x_c),
    .io_y_ppn(tlb_ppn_data_barrier_4_io_y_ppn),
    .io_y_u(tlb_ppn_data_barrier_4_io_y_u),
    .io_y_ae(tlb_ppn_data_barrier_4_io_y_ae),
    .io_y_sw(tlb_ppn_data_barrier_4_io_y_sw),
    .io_y_sx(tlb_ppn_data_barrier_4_io_y_sx),
    .io_y_sr(tlb_ppn_data_barrier_4_io_y_sr),
    .io_y_pw(tlb_ppn_data_barrier_4_io_y_pw),
    .io_y_px(tlb_ppn_data_barrier_4_io_y_px),
    .io_y_pr(tlb_ppn_data_barrier_4_io_y_pr),
    .io_y_ppp(tlb_ppn_data_barrier_4_io_y_ppp),
    .io_y_pal(tlb_ppn_data_barrier_4_io_y_pal),
    .io_y_paa(tlb_ppn_data_barrier_4_io_y_paa),
    .io_y_eff(tlb_ppn_data_barrier_4_io_y_eff),
    .io_y_c(tlb_ppn_data_barrier_4_io_y_c)
  );
  OptimizationBarrier tlb_ppn_data_barrier_5 ( // @[package.scala 236:25]
    .io_x_ppn(tlb_ppn_data_barrier_5_io_x_ppn),
    .io_x_u(tlb_ppn_data_barrier_5_io_x_u),
    .io_x_ae(tlb_ppn_data_barrier_5_io_x_ae),
    .io_x_sw(tlb_ppn_data_barrier_5_io_x_sw),
    .io_x_sx(tlb_ppn_data_barrier_5_io_x_sx),
    .io_x_sr(tlb_ppn_data_barrier_5_io_x_sr),
    .io_x_pw(tlb_ppn_data_barrier_5_io_x_pw),
    .io_x_px(tlb_ppn_data_barrier_5_io_x_px),
    .io_x_pr(tlb_ppn_data_barrier_5_io_x_pr),
    .io_x_ppp(tlb_ppn_data_barrier_5_io_x_ppp),
    .io_x_pal(tlb_ppn_data_barrier_5_io_x_pal),
    .io_x_paa(tlb_ppn_data_barrier_5_io_x_paa),
    .io_x_eff(tlb_ppn_data_barrier_5_io_x_eff),
    .io_x_c(tlb_ppn_data_barrier_5_io_x_c),
    .io_y_ppn(tlb_ppn_data_barrier_5_io_y_ppn),
    .io_y_u(tlb_ppn_data_barrier_5_io_y_u),
    .io_y_ae(tlb_ppn_data_barrier_5_io_y_ae),
    .io_y_sw(tlb_ppn_data_barrier_5_io_y_sw),
    .io_y_sx(tlb_ppn_data_barrier_5_io_y_sx),
    .io_y_sr(tlb_ppn_data_barrier_5_io_y_sr),
    .io_y_pw(tlb_ppn_data_barrier_5_io_y_pw),
    .io_y_px(tlb_ppn_data_barrier_5_io_y_px),
    .io_y_pr(tlb_ppn_data_barrier_5_io_y_pr),
    .io_y_ppp(tlb_ppn_data_barrier_5_io_y_ppp),
    .io_y_pal(tlb_ppn_data_barrier_5_io_y_pal),
    .io_y_paa(tlb_ppn_data_barrier_5_io_y_paa),
    .io_y_eff(tlb_ppn_data_barrier_5_io_y_eff),
    .io_y_c(tlb_ppn_data_barrier_5_io_y_c)
  );
  OptimizationBarrier tlb_ppn_data_barrier_6 ( // @[package.scala 236:25]
    .io_x_ppn(tlb_ppn_data_barrier_6_io_x_ppn),
    .io_x_u(tlb_ppn_data_barrier_6_io_x_u),
    .io_x_ae(tlb_ppn_data_barrier_6_io_x_ae),
    .io_x_sw(tlb_ppn_data_barrier_6_io_x_sw),
    .io_x_sx(tlb_ppn_data_barrier_6_io_x_sx),
    .io_x_sr(tlb_ppn_data_barrier_6_io_x_sr),
    .io_x_pw(tlb_ppn_data_barrier_6_io_x_pw),
    .io_x_px(tlb_ppn_data_barrier_6_io_x_px),
    .io_x_pr(tlb_ppn_data_barrier_6_io_x_pr),
    .io_x_ppp(tlb_ppn_data_barrier_6_io_x_ppp),
    .io_x_pal(tlb_ppn_data_barrier_6_io_x_pal),
    .io_x_paa(tlb_ppn_data_barrier_6_io_x_paa),
    .io_x_eff(tlb_ppn_data_barrier_6_io_x_eff),
    .io_x_c(tlb_ppn_data_barrier_6_io_x_c),
    .io_y_ppn(tlb_ppn_data_barrier_6_io_y_ppn),
    .io_y_u(tlb_ppn_data_barrier_6_io_y_u),
    .io_y_ae(tlb_ppn_data_barrier_6_io_y_ae),
    .io_y_sw(tlb_ppn_data_barrier_6_io_y_sw),
    .io_y_sx(tlb_ppn_data_barrier_6_io_y_sx),
    .io_y_sr(tlb_ppn_data_barrier_6_io_y_sr),
    .io_y_pw(tlb_ppn_data_barrier_6_io_y_pw),
    .io_y_px(tlb_ppn_data_barrier_6_io_y_px),
    .io_y_pr(tlb_ppn_data_barrier_6_io_y_pr),
    .io_y_ppp(tlb_ppn_data_barrier_6_io_y_ppp),
    .io_y_pal(tlb_ppn_data_barrier_6_io_y_pal),
    .io_y_paa(tlb_ppn_data_barrier_6_io_y_paa),
    .io_y_eff(tlb_ppn_data_barrier_6_io_y_eff),
    .io_y_c(tlb_ppn_data_barrier_6_io_y_c)
  );
  OptimizationBarrier tlb_ppn_data_barrier_7 ( // @[package.scala 236:25]
    .io_x_ppn(tlb_ppn_data_barrier_7_io_x_ppn),
    .io_x_u(tlb_ppn_data_barrier_7_io_x_u),
    .io_x_ae(tlb_ppn_data_barrier_7_io_x_ae),
    .io_x_sw(tlb_ppn_data_barrier_7_io_x_sw),
    .io_x_sx(tlb_ppn_data_barrier_7_io_x_sx),
    .io_x_sr(tlb_ppn_data_barrier_7_io_x_sr),
    .io_x_pw(tlb_ppn_data_barrier_7_io_x_pw),
    .io_x_px(tlb_ppn_data_barrier_7_io_x_px),
    .io_x_pr(tlb_ppn_data_barrier_7_io_x_pr),
    .io_x_ppp(tlb_ppn_data_barrier_7_io_x_ppp),
    .io_x_pal(tlb_ppn_data_barrier_7_io_x_pal),
    .io_x_paa(tlb_ppn_data_barrier_7_io_x_paa),
    .io_x_eff(tlb_ppn_data_barrier_7_io_x_eff),
    .io_x_c(tlb_ppn_data_barrier_7_io_x_c),
    .io_y_ppn(tlb_ppn_data_barrier_7_io_y_ppn),
    .io_y_u(tlb_ppn_data_barrier_7_io_y_u),
    .io_y_ae(tlb_ppn_data_barrier_7_io_y_ae),
    .io_y_sw(tlb_ppn_data_barrier_7_io_y_sw),
    .io_y_sx(tlb_ppn_data_barrier_7_io_y_sx),
    .io_y_sr(tlb_ppn_data_barrier_7_io_y_sr),
    .io_y_pw(tlb_ppn_data_barrier_7_io_y_pw),
    .io_y_px(tlb_ppn_data_barrier_7_io_y_px),
    .io_y_pr(tlb_ppn_data_barrier_7_io_y_pr),
    .io_y_ppp(tlb_ppn_data_barrier_7_io_y_ppp),
    .io_y_pal(tlb_ppn_data_barrier_7_io_y_pal),
    .io_y_paa(tlb_ppn_data_barrier_7_io_y_paa),
    .io_y_eff(tlb_ppn_data_barrier_7_io_y_eff),
    .io_y_c(tlb_ppn_data_barrier_7_io_y_c)
  );
  OptimizationBarrier tlb_ppn_data_barrier_8 ( // @[package.scala 236:25]
    .io_x_ppn(tlb_ppn_data_barrier_8_io_x_ppn),
    .io_x_u(tlb_ppn_data_barrier_8_io_x_u),
    .io_x_ae(tlb_ppn_data_barrier_8_io_x_ae),
    .io_x_sw(tlb_ppn_data_barrier_8_io_x_sw),
    .io_x_sx(tlb_ppn_data_barrier_8_io_x_sx),
    .io_x_sr(tlb_ppn_data_barrier_8_io_x_sr),
    .io_x_pw(tlb_ppn_data_barrier_8_io_x_pw),
    .io_x_px(tlb_ppn_data_barrier_8_io_x_px),
    .io_x_pr(tlb_ppn_data_barrier_8_io_x_pr),
    .io_x_ppp(tlb_ppn_data_barrier_8_io_x_ppp),
    .io_x_pal(tlb_ppn_data_barrier_8_io_x_pal),
    .io_x_paa(tlb_ppn_data_barrier_8_io_x_paa),
    .io_x_eff(tlb_ppn_data_barrier_8_io_x_eff),
    .io_x_c(tlb_ppn_data_barrier_8_io_x_c),
    .io_y_ppn(tlb_ppn_data_barrier_8_io_y_ppn),
    .io_y_u(tlb_ppn_data_barrier_8_io_y_u),
    .io_y_ae(tlb_ppn_data_barrier_8_io_y_ae),
    .io_y_sw(tlb_ppn_data_barrier_8_io_y_sw),
    .io_y_sx(tlb_ppn_data_barrier_8_io_y_sx),
    .io_y_sr(tlb_ppn_data_barrier_8_io_y_sr),
    .io_y_pw(tlb_ppn_data_barrier_8_io_y_pw),
    .io_y_px(tlb_ppn_data_barrier_8_io_y_px),
    .io_y_pr(tlb_ppn_data_barrier_8_io_y_pr),
    .io_y_ppp(tlb_ppn_data_barrier_8_io_y_ppp),
    .io_y_pal(tlb_ppn_data_barrier_8_io_y_pal),
    .io_y_paa(tlb_ppn_data_barrier_8_io_y_paa),
    .io_y_eff(tlb_ppn_data_barrier_8_io_y_eff),
    .io_y_c(tlb_ppn_data_barrier_8_io_y_c)
  );
  OptimizationBarrier tlb_ppn_data_barrier_9 ( // @[package.scala 236:25]
    .io_x_ppn(tlb_ppn_data_barrier_9_io_x_ppn),
    .io_x_u(tlb_ppn_data_barrier_9_io_x_u),
    .io_x_ae(tlb_ppn_data_barrier_9_io_x_ae),
    .io_x_sw(tlb_ppn_data_barrier_9_io_x_sw),
    .io_x_sx(tlb_ppn_data_barrier_9_io_x_sx),
    .io_x_sr(tlb_ppn_data_barrier_9_io_x_sr),
    .io_x_pw(tlb_ppn_data_barrier_9_io_x_pw),
    .io_x_px(tlb_ppn_data_barrier_9_io_x_px),
    .io_x_pr(tlb_ppn_data_barrier_9_io_x_pr),
    .io_x_ppp(tlb_ppn_data_barrier_9_io_x_ppp),
    .io_x_pal(tlb_ppn_data_barrier_9_io_x_pal),
    .io_x_paa(tlb_ppn_data_barrier_9_io_x_paa),
    .io_x_eff(tlb_ppn_data_barrier_9_io_x_eff),
    .io_x_c(tlb_ppn_data_barrier_9_io_x_c),
    .io_y_ppn(tlb_ppn_data_barrier_9_io_y_ppn),
    .io_y_u(tlb_ppn_data_barrier_9_io_y_u),
    .io_y_ae(tlb_ppn_data_barrier_9_io_y_ae),
    .io_y_sw(tlb_ppn_data_barrier_9_io_y_sw),
    .io_y_sx(tlb_ppn_data_barrier_9_io_y_sx),
    .io_y_sr(tlb_ppn_data_barrier_9_io_y_sr),
    .io_y_pw(tlb_ppn_data_barrier_9_io_y_pw),
    .io_y_px(tlb_ppn_data_barrier_9_io_y_px),
    .io_y_pr(tlb_ppn_data_barrier_9_io_y_pr),
    .io_y_ppp(tlb_ppn_data_barrier_9_io_y_ppp),
    .io_y_pal(tlb_ppn_data_barrier_9_io_y_pal),
    .io_y_paa(tlb_ppn_data_barrier_9_io_y_paa),
    .io_y_eff(tlb_ppn_data_barrier_9_io_y_eff),
    .io_y_c(tlb_ppn_data_barrier_9_io_y_c)
  );
  OptimizationBarrier tlb_ppn_data_barrier_10 ( // @[package.scala 236:25]
    .io_x_ppn(tlb_ppn_data_barrier_10_io_x_ppn),
    .io_x_u(tlb_ppn_data_barrier_10_io_x_u),
    .io_x_ae(tlb_ppn_data_barrier_10_io_x_ae),
    .io_x_sw(tlb_ppn_data_barrier_10_io_x_sw),
    .io_x_sx(tlb_ppn_data_barrier_10_io_x_sx),
    .io_x_sr(tlb_ppn_data_barrier_10_io_x_sr),
    .io_x_pw(tlb_ppn_data_barrier_10_io_x_pw),
    .io_x_px(tlb_ppn_data_barrier_10_io_x_px),
    .io_x_pr(tlb_ppn_data_barrier_10_io_x_pr),
    .io_x_ppp(tlb_ppn_data_barrier_10_io_x_ppp),
    .io_x_pal(tlb_ppn_data_barrier_10_io_x_pal),
    .io_x_paa(tlb_ppn_data_barrier_10_io_x_paa),
    .io_x_eff(tlb_ppn_data_barrier_10_io_x_eff),
    .io_x_c(tlb_ppn_data_barrier_10_io_x_c),
    .io_y_ppn(tlb_ppn_data_barrier_10_io_y_ppn),
    .io_y_u(tlb_ppn_data_barrier_10_io_y_u),
    .io_y_ae(tlb_ppn_data_barrier_10_io_y_ae),
    .io_y_sw(tlb_ppn_data_barrier_10_io_y_sw),
    .io_y_sx(tlb_ppn_data_barrier_10_io_y_sx),
    .io_y_sr(tlb_ppn_data_barrier_10_io_y_sr),
    .io_y_pw(tlb_ppn_data_barrier_10_io_y_pw),
    .io_y_px(tlb_ppn_data_barrier_10_io_y_px),
    .io_y_pr(tlb_ppn_data_barrier_10_io_y_pr),
    .io_y_ppp(tlb_ppn_data_barrier_10_io_y_ppp),
    .io_y_pal(tlb_ppn_data_barrier_10_io_y_pal),
    .io_y_paa(tlb_ppn_data_barrier_10_io_y_paa),
    .io_y_eff(tlb_ppn_data_barrier_10_io_y_eff),
    .io_y_c(tlb_ppn_data_barrier_10_io_y_c)
  );
  OptimizationBarrier tlb_ppn_data_barrier_11 ( // @[package.scala 236:25]
    .io_x_ppn(tlb_ppn_data_barrier_11_io_x_ppn),
    .io_x_u(tlb_ppn_data_barrier_11_io_x_u),
    .io_x_ae(tlb_ppn_data_barrier_11_io_x_ae),
    .io_x_sw(tlb_ppn_data_barrier_11_io_x_sw),
    .io_x_sx(tlb_ppn_data_barrier_11_io_x_sx),
    .io_x_sr(tlb_ppn_data_barrier_11_io_x_sr),
    .io_x_pw(tlb_ppn_data_barrier_11_io_x_pw),
    .io_x_px(tlb_ppn_data_barrier_11_io_x_px),
    .io_x_pr(tlb_ppn_data_barrier_11_io_x_pr),
    .io_x_ppp(tlb_ppn_data_barrier_11_io_x_ppp),
    .io_x_pal(tlb_ppn_data_barrier_11_io_x_pal),
    .io_x_paa(tlb_ppn_data_barrier_11_io_x_paa),
    .io_x_eff(tlb_ppn_data_barrier_11_io_x_eff),
    .io_x_c(tlb_ppn_data_barrier_11_io_x_c),
    .io_y_ppn(tlb_ppn_data_barrier_11_io_y_ppn),
    .io_y_u(tlb_ppn_data_barrier_11_io_y_u),
    .io_y_ae(tlb_ppn_data_barrier_11_io_y_ae),
    .io_y_sw(tlb_ppn_data_barrier_11_io_y_sw),
    .io_y_sx(tlb_ppn_data_barrier_11_io_y_sx),
    .io_y_sr(tlb_ppn_data_barrier_11_io_y_sr),
    .io_y_pw(tlb_ppn_data_barrier_11_io_y_pw),
    .io_y_px(tlb_ppn_data_barrier_11_io_y_px),
    .io_y_pr(tlb_ppn_data_barrier_11_io_y_pr),
    .io_y_ppp(tlb_ppn_data_barrier_11_io_y_ppp),
    .io_y_pal(tlb_ppn_data_barrier_11_io_y_pal),
    .io_y_paa(tlb_ppn_data_barrier_11_io_y_paa),
    .io_y_eff(tlb_ppn_data_barrier_11_io_y_eff),
    .io_y_c(tlb_ppn_data_barrier_11_io_y_c)
  );
  OptimizationBarrier tlb_ppn_data_barrier_12 ( // @[package.scala 236:25]
    .io_x_ppn(tlb_ppn_data_barrier_12_io_x_ppn),
    .io_x_u(tlb_ppn_data_barrier_12_io_x_u),
    .io_x_ae(tlb_ppn_data_barrier_12_io_x_ae),
    .io_x_sw(tlb_ppn_data_barrier_12_io_x_sw),
    .io_x_sx(tlb_ppn_data_barrier_12_io_x_sx),
    .io_x_sr(tlb_ppn_data_barrier_12_io_x_sr),
    .io_x_pw(tlb_ppn_data_barrier_12_io_x_pw),
    .io_x_px(tlb_ppn_data_barrier_12_io_x_px),
    .io_x_pr(tlb_ppn_data_barrier_12_io_x_pr),
    .io_x_ppp(tlb_ppn_data_barrier_12_io_x_ppp),
    .io_x_pal(tlb_ppn_data_barrier_12_io_x_pal),
    .io_x_paa(tlb_ppn_data_barrier_12_io_x_paa),
    .io_x_eff(tlb_ppn_data_barrier_12_io_x_eff),
    .io_x_c(tlb_ppn_data_barrier_12_io_x_c),
    .io_y_ppn(tlb_ppn_data_barrier_12_io_y_ppn),
    .io_y_u(tlb_ppn_data_barrier_12_io_y_u),
    .io_y_ae(tlb_ppn_data_barrier_12_io_y_ae),
    .io_y_sw(tlb_ppn_data_barrier_12_io_y_sw),
    .io_y_sx(tlb_ppn_data_barrier_12_io_y_sx),
    .io_y_sr(tlb_ppn_data_barrier_12_io_y_sr),
    .io_y_pw(tlb_ppn_data_barrier_12_io_y_pw),
    .io_y_px(tlb_ppn_data_barrier_12_io_y_px),
    .io_y_pr(tlb_ppn_data_barrier_12_io_y_pr),
    .io_y_ppp(tlb_ppn_data_barrier_12_io_y_ppp),
    .io_y_pal(tlb_ppn_data_barrier_12_io_y_pal),
    .io_y_paa(tlb_ppn_data_barrier_12_io_y_paa),
    .io_y_eff(tlb_ppn_data_barrier_12_io_y_eff),
    .io_y_c(tlb_ppn_data_barrier_12_io_y_c)
  );
  OptimizationBarrier tlb_entries_barrier ( // @[package.scala 236:25]
    .io_x_ppn(tlb_entries_barrier_io_x_ppn),
    .io_x_u(tlb_entries_barrier_io_x_u),
    .io_x_ae(tlb_entries_barrier_io_x_ae),
    .io_x_sw(tlb_entries_barrier_io_x_sw),
    .io_x_sx(tlb_entries_barrier_io_x_sx),
    .io_x_sr(tlb_entries_barrier_io_x_sr),
    .io_x_pw(tlb_entries_barrier_io_x_pw),
    .io_x_px(tlb_entries_barrier_io_x_px),
    .io_x_pr(tlb_entries_barrier_io_x_pr),
    .io_x_ppp(tlb_entries_barrier_io_x_ppp),
    .io_x_pal(tlb_entries_barrier_io_x_pal),
    .io_x_paa(tlb_entries_barrier_io_x_paa),
    .io_x_eff(tlb_entries_barrier_io_x_eff),
    .io_x_c(tlb_entries_barrier_io_x_c),
    .io_y_ppn(tlb_entries_barrier_io_y_ppn),
    .io_y_u(tlb_entries_barrier_io_y_u),
    .io_y_ae(tlb_entries_barrier_io_y_ae),
    .io_y_sw(tlb_entries_barrier_io_y_sw),
    .io_y_sx(tlb_entries_barrier_io_y_sx),
    .io_y_sr(tlb_entries_barrier_io_y_sr),
    .io_y_pw(tlb_entries_barrier_io_y_pw),
    .io_y_px(tlb_entries_barrier_io_y_px),
    .io_y_pr(tlb_entries_barrier_io_y_pr),
    .io_y_ppp(tlb_entries_barrier_io_y_ppp),
    .io_y_pal(tlb_entries_barrier_io_y_pal),
    .io_y_paa(tlb_entries_barrier_io_y_paa),
    .io_y_eff(tlb_entries_barrier_io_y_eff),
    .io_y_c(tlb_entries_barrier_io_y_c)
  );
  OptimizationBarrier tlb_entries_barrier_1 ( // @[package.scala 236:25]
    .io_x_ppn(tlb_entries_barrier_1_io_x_ppn),
    .io_x_u(tlb_entries_barrier_1_io_x_u),
    .io_x_ae(tlb_entries_barrier_1_io_x_ae),
    .io_x_sw(tlb_entries_barrier_1_io_x_sw),
    .io_x_sx(tlb_entries_barrier_1_io_x_sx),
    .io_x_sr(tlb_entries_barrier_1_io_x_sr),
    .io_x_pw(tlb_entries_barrier_1_io_x_pw),
    .io_x_px(tlb_entries_barrier_1_io_x_px),
    .io_x_pr(tlb_entries_barrier_1_io_x_pr),
    .io_x_ppp(tlb_entries_barrier_1_io_x_ppp),
    .io_x_pal(tlb_entries_barrier_1_io_x_pal),
    .io_x_paa(tlb_entries_barrier_1_io_x_paa),
    .io_x_eff(tlb_entries_barrier_1_io_x_eff),
    .io_x_c(tlb_entries_barrier_1_io_x_c),
    .io_y_ppn(tlb_entries_barrier_1_io_y_ppn),
    .io_y_u(tlb_entries_barrier_1_io_y_u),
    .io_y_ae(tlb_entries_barrier_1_io_y_ae),
    .io_y_sw(tlb_entries_barrier_1_io_y_sw),
    .io_y_sx(tlb_entries_barrier_1_io_y_sx),
    .io_y_sr(tlb_entries_barrier_1_io_y_sr),
    .io_y_pw(tlb_entries_barrier_1_io_y_pw),
    .io_y_px(tlb_entries_barrier_1_io_y_px),
    .io_y_pr(tlb_entries_barrier_1_io_y_pr),
    .io_y_ppp(tlb_entries_barrier_1_io_y_ppp),
    .io_y_pal(tlb_entries_barrier_1_io_y_pal),
    .io_y_paa(tlb_entries_barrier_1_io_y_paa),
    .io_y_eff(tlb_entries_barrier_1_io_y_eff),
    .io_y_c(tlb_entries_barrier_1_io_y_c)
  );
  OptimizationBarrier tlb_entries_barrier_2 ( // @[package.scala 236:25]
    .io_x_ppn(tlb_entries_barrier_2_io_x_ppn),
    .io_x_u(tlb_entries_barrier_2_io_x_u),
    .io_x_ae(tlb_entries_barrier_2_io_x_ae),
    .io_x_sw(tlb_entries_barrier_2_io_x_sw),
    .io_x_sx(tlb_entries_barrier_2_io_x_sx),
    .io_x_sr(tlb_entries_barrier_2_io_x_sr),
    .io_x_pw(tlb_entries_barrier_2_io_x_pw),
    .io_x_px(tlb_entries_barrier_2_io_x_px),
    .io_x_pr(tlb_entries_barrier_2_io_x_pr),
    .io_x_ppp(tlb_entries_barrier_2_io_x_ppp),
    .io_x_pal(tlb_entries_barrier_2_io_x_pal),
    .io_x_paa(tlb_entries_barrier_2_io_x_paa),
    .io_x_eff(tlb_entries_barrier_2_io_x_eff),
    .io_x_c(tlb_entries_barrier_2_io_x_c),
    .io_y_ppn(tlb_entries_barrier_2_io_y_ppn),
    .io_y_u(tlb_entries_barrier_2_io_y_u),
    .io_y_ae(tlb_entries_barrier_2_io_y_ae),
    .io_y_sw(tlb_entries_barrier_2_io_y_sw),
    .io_y_sx(tlb_entries_barrier_2_io_y_sx),
    .io_y_sr(tlb_entries_barrier_2_io_y_sr),
    .io_y_pw(tlb_entries_barrier_2_io_y_pw),
    .io_y_px(tlb_entries_barrier_2_io_y_px),
    .io_y_pr(tlb_entries_barrier_2_io_y_pr),
    .io_y_ppp(tlb_entries_barrier_2_io_y_ppp),
    .io_y_pal(tlb_entries_barrier_2_io_y_pal),
    .io_y_paa(tlb_entries_barrier_2_io_y_paa),
    .io_y_eff(tlb_entries_barrier_2_io_y_eff),
    .io_y_c(tlb_entries_barrier_2_io_y_c)
  );
  OptimizationBarrier tlb_entries_barrier_3 ( // @[package.scala 236:25]
    .io_x_ppn(tlb_entries_barrier_3_io_x_ppn),
    .io_x_u(tlb_entries_barrier_3_io_x_u),
    .io_x_ae(tlb_entries_barrier_3_io_x_ae),
    .io_x_sw(tlb_entries_barrier_3_io_x_sw),
    .io_x_sx(tlb_entries_barrier_3_io_x_sx),
    .io_x_sr(tlb_entries_barrier_3_io_x_sr),
    .io_x_pw(tlb_entries_barrier_3_io_x_pw),
    .io_x_px(tlb_entries_barrier_3_io_x_px),
    .io_x_pr(tlb_entries_barrier_3_io_x_pr),
    .io_x_ppp(tlb_entries_barrier_3_io_x_ppp),
    .io_x_pal(tlb_entries_barrier_3_io_x_pal),
    .io_x_paa(tlb_entries_barrier_3_io_x_paa),
    .io_x_eff(tlb_entries_barrier_3_io_x_eff),
    .io_x_c(tlb_entries_barrier_3_io_x_c),
    .io_y_ppn(tlb_entries_barrier_3_io_y_ppn),
    .io_y_u(tlb_entries_barrier_3_io_y_u),
    .io_y_ae(tlb_entries_barrier_3_io_y_ae),
    .io_y_sw(tlb_entries_barrier_3_io_y_sw),
    .io_y_sx(tlb_entries_barrier_3_io_y_sx),
    .io_y_sr(tlb_entries_barrier_3_io_y_sr),
    .io_y_pw(tlb_entries_barrier_3_io_y_pw),
    .io_y_px(tlb_entries_barrier_3_io_y_px),
    .io_y_pr(tlb_entries_barrier_3_io_y_pr),
    .io_y_ppp(tlb_entries_barrier_3_io_y_ppp),
    .io_y_pal(tlb_entries_barrier_3_io_y_pal),
    .io_y_paa(tlb_entries_barrier_3_io_y_paa),
    .io_y_eff(tlb_entries_barrier_3_io_y_eff),
    .io_y_c(tlb_entries_barrier_3_io_y_c)
  );
  OptimizationBarrier tlb_entries_barrier_4 ( // @[package.scala 236:25]
    .io_x_ppn(tlb_entries_barrier_4_io_x_ppn),
    .io_x_u(tlb_entries_barrier_4_io_x_u),
    .io_x_ae(tlb_entries_barrier_4_io_x_ae),
    .io_x_sw(tlb_entries_barrier_4_io_x_sw),
    .io_x_sx(tlb_entries_barrier_4_io_x_sx),
    .io_x_sr(tlb_entries_barrier_4_io_x_sr),
    .io_x_pw(tlb_entries_barrier_4_io_x_pw),
    .io_x_px(tlb_entries_barrier_4_io_x_px),
    .io_x_pr(tlb_entries_barrier_4_io_x_pr),
    .io_x_ppp(tlb_entries_barrier_4_io_x_ppp),
    .io_x_pal(tlb_entries_barrier_4_io_x_pal),
    .io_x_paa(tlb_entries_barrier_4_io_x_paa),
    .io_x_eff(tlb_entries_barrier_4_io_x_eff),
    .io_x_c(tlb_entries_barrier_4_io_x_c),
    .io_y_ppn(tlb_entries_barrier_4_io_y_ppn),
    .io_y_u(tlb_entries_barrier_4_io_y_u),
    .io_y_ae(tlb_entries_barrier_4_io_y_ae),
    .io_y_sw(tlb_entries_barrier_4_io_y_sw),
    .io_y_sx(tlb_entries_barrier_4_io_y_sx),
    .io_y_sr(tlb_entries_barrier_4_io_y_sr),
    .io_y_pw(tlb_entries_barrier_4_io_y_pw),
    .io_y_px(tlb_entries_barrier_4_io_y_px),
    .io_y_pr(tlb_entries_barrier_4_io_y_pr),
    .io_y_ppp(tlb_entries_barrier_4_io_y_ppp),
    .io_y_pal(tlb_entries_barrier_4_io_y_pal),
    .io_y_paa(tlb_entries_barrier_4_io_y_paa),
    .io_y_eff(tlb_entries_barrier_4_io_y_eff),
    .io_y_c(tlb_entries_barrier_4_io_y_c)
  );
  OptimizationBarrier tlb_entries_barrier_5 ( // @[package.scala 236:25]
    .io_x_ppn(tlb_entries_barrier_5_io_x_ppn),
    .io_x_u(tlb_entries_barrier_5_io_x_u),
    .io_x_ae(tlb_entries_barrier_5_io_x_ae),
    .io_x_sw(tlb_entries_barrier_5_io_x_sw),
    .io_x_sx(tlb_entries_barrier_5_io_x_sx),
    .io_x_sr(tlb_entries_barrier_5_io_x_sr),
    .io_x_pw(tlb_entries_barrier_5_io_x_pw),
    .io_x_px(tlb_entries_barrier_5_io_x_px),
    .io_x_pr(tlb_entries_barrier_5_io_x_pr),
    .io_x_ppp(tlb_entries_barrier_5_io_x_ppp),
    .io_x_pal(tlb_entries_barrier_5_io_x_pal),
    .io_x_paa(tlb_entries_barrier_5_io_x_paa),
    .io_x_eff(tlb_entries_barrier_5_io_x_eff),
    .io_x_c(tlb_entries_barrier_5_io_x_c),
    .io_y_ppn(tlb_entries_barrier_5_io_y_ppn),
    .io_y_u(tlb_entries_barrier_5_io_y_u),
    .io_y_ae(tlb_entries_barrier_5_io_y_ae),
    .io_y_sw(tlb_entries_barrier_5_io_y_sw),
    .io_y_sx(tlb_entries_barrier_5_io_y_sx),
    .io_y_sr(tlb_entries_barrier_5_io_y_sr),
    .io_y_pw(tlb_entries_barrier_5_io_y_pw),
    .io_y_px(tlb_entries_barrier_5_io_y_px),
    .io_y_pr(tlb_entries_barrier_5_io_y_pr),
    .io_y_ppp(tlb_entries_barrier_5_io_y_ppp),
    .io_y_pal(tlb_entries_barrier_5_io_y_pal),
    .io_y_paa(tlb_entries_barrier_5_io_y_paa),
    .io_y_eff(tlb_entries_barrier_5_io_y_eff),
    .io_y_c(tlb_entries_barrier_5_io_y_c)
  );
  OptimizationBarrier tlb_entries_barrier_6 ( // @[package.scala 236:25]
    .io_x_ppn(tlb_entries_barrier_6_io_x_ppn),
    .io_x_u(tlb_entries_barrier_6_io_x_u),
    .io_x_ae(tlb_entries_barrier_6_io_x_ae),
    .io_x_sw(tlb_entries_barrier_6_io_x_sw),
    .io_x_sx(tlb_entries_barrier_6_io_x_sx),
    .io_x_sr(tlb_entries_barrier_6_io_x_sr),
    .io_x_pw(tlb_entries_barrier_6_io_x_pw),
    .io_x_px(tlb_entries_barrier_6_io_x_px),
    .io_x_pr(tlb_entries_barrier_6_io_x_pr),
    .io_x_ppp(tlb_entries_barrier_6_io_x_ppp),
    .io_x_pal(tlb_entries_barrier_6_io_x_pal),
    .io_x_paa(tlb_entries_barrier_6_io_x_paa),
    .io_x_eff(tlb_entries_barrier_6_io_x_eff),
    .io_x_c(tlb_entries_barrier_6_io_x_c),
    .io_y_ppn(tlb_entries_barrier_6_io_y_ppn),
    .io_y_u(tlb_entries_barrier_6_io_y_u),
    .io_y_ae(tlb_entries_barrier_6_io_y_ae),
    .io_y_sw(tlb_entries_barrier_6_io_y_sw),
    .io_y_sx(tlb_entries_barrier_6_io_y_sx),
    .io_y_sr(tlb_entries_barrier_6_io_y_sr),
    .io_y_pw(tlb_entries_barrier_6_io_y_pw),
    .io_y_px(tlb_entries_barrier_6_io_y_px),
    .io_y_pr(tlb_entries_barrier_6_io_y_pr),
    .io_y_ppp(tlb_entries_barrier_6_io_y_ppp),
    .io_y_pal(tlb_entries_barrier_6_io_y_pal),
    .io_y_paa(tlb_entries_barrier_6_io_y_paa),
    .io_y_eff(tlb_entries_barrier_6_io_y_eff),
    .io_y_c(tlb_entries_barrier_6_io_y_c)
  );
  OptimizationBarrier tlb_entries_barrier_7 ( // @[package.scala 236:25]
    .io_x_ppn(tlb_entries_barrier_7_io_x_ppn),
    .io_x_u(tlb_entries_barrier_7_io_x_u),
    .io_x_ae(tlb_entries_barrier_7_io_x_ae),
    .io_x_sw(tlb_entries_barrier_7_io_x_sw),
    .io_x_sx(tlb_entries_barrier_7_io_x_sx),
    .io_x_sr(tlb_entries_barrier_7_io_x_sr),
    .io_x_pw(tlb_entries_barrier_7_io_x_pw),
    .io_x_px(tlb_entries_barrier_7_io_x_px),
    .io_x_pr(tlb_entries_barrier_7_io_x_pr),
    .io_x_ppp(tlb_entries_barrier_7_io_x_ppp),
    .io_x_pal(tlb_entries_barrier_7_io_x_pal),
    .io_x_paa(tlb_entries_barrier_7_io_x_paa),
    .io_x_eff(tlb_entries_barrier_7_io_x_eff),
    .io_x_c(tlb_entries_barrier_7_io_x_c),
    .io_y_ppn(tlb_entries_barrier_7_io_y_ppn),
    .io_y_u(tlb_entries_barrier_7_io_y_u),
    .io_y_ae(tlb_entries_barrier_7_io_y_ae),
    .io_y_sw(tlb_entries_barrier_7_io_y_sw),
    .io_y_sx(tlb_entries_barrier_7_io_y_sx),
    .io_y_sr(tlb_entries_barrier_7_io_y_sr),
    .io_y_pw(tlb_entries_barrier_7_io_y_pw),
    .io_y_px(tlb_entries_barrier_7_io_y_px),
    .io_y_pr(tlb_entries_barrier_7_io_y_pr),
    .io_y_ppp(tlb_entries_barrier_7_io_y_ppp),
    .io_y_pal(tlb_entries_barrier_7_io_y_pal),
    .io_y_paa(tlb_entries_barrier_7_io_y_paa),
    .io_y_eff(tlb_entries_barrier_7_io_y_eff),
    .io_y_c(tlb_entries_barrier_7_io_y_c)
  );
  OptimizationBarrier tlb_entries_barrier_8 ( // @[package.scala 236:25]
    .io_x_ppn(tlb_entries_barrier_8_io_x_ppn),
    .io_x_u(tlb_entries_barrier_8_io_x_u),
    .io_x_ae(tlb_entries_barrier_8_io_x_ae),
    .io_x_sw(tlb_entries_barrier_8_io_x_sw),
    .io_x_sx(tlb_entries_barrier_8_io_x_sx),
    .io_x_sr(tlb_entries_barrier_8_io_x_sr),
    .io_x_pw(tlb_entries_barrier_8_io_x_pw),
    .io_x_px(tlb_entries_barrier_8_io_x_px),
    .io_x_pr(tlb_entries_barrier_8_io_x_pr),
    .io_x_ppp(tlb_entries_barrier_8_io_x_ppp),
    .io_x_pal(tlb_entries_barrier_8_io_x_pal),
    .io_x_paa(tlb_entries_barrier_8_io_x_paa),
    .io_x_eff(tlb_entries_barrier_8_io_x_eff),
    .io_x_c(tlb_entries_barrier_8_io_x_c),
    .io_y_ppn(tlb_entries_barrier_8_io_y_ppn),
    .io_y_u(tlb_entries_barrier_8_io_y_u),
    .io_y_ae(tlb_entries_barrier_8_io_y_ae),
    .io_y_sw(tlb_entries_barrier_8_io_y_sw),
    .io_y_sx(tlb_entries_barrier_8_io_y_sx),
    .io_y_sr(tlb_entries_barrier_8_io_y_sr),
    .io_y_pw(tlb_entries_barrier_8_io_y_pw),
    .io_y_px(tlb_entries_barrier_8_io_y_px),
    .io_y_pr(tlb_entries_barrier_8_io_y_pr),
    .io_y_ppp(tlb_entries_barrier_8_io_y_ppp),
    .io_y_pal(tlb_entries_barrier_8_io_y_pal),
    .io_y_paa(tlb_entries_barrier_8_io_y_paa),
    .io_y_eff(tlb_entries_barrier_8_io_y_eff),
    .io_y_c(tlb_entries_barrier_8_io_y_c)
  );
  OptimizationBarrier tlb_entries_barrier_9 ( // @[package.scala 236:25]
    .io_x_ppn(tlb_entries_barrier_9_io_x_ppn),
    .io_x_u(tlb_entries_barrier_9_io_x_u),
    .io_x_ae(tlb_entries_barrier_9_io_x_ae),
    .io_x_sw(tlb_entries_barrier_9_io_x_sw),
    .io_x_sx(tlb_entries_barrier_9_io_x_sx),
    .io_x_sr(tlb_entries_barrier_9_io_x_sr),
    .io_x_pw(tlb_entries_barrier_9_io_x_pw),
    .io_x_px(tlb_entries_barrier_9_io_x_px),
    .io_x_pr(tlb_entries_barrier_9_io_x_pr),
    .io_x_ppp(tlb_entries_barrier_9_io_x_ppp),
    .io_x_pal(tlb_entries_barrier_9_io_x_pal),
    .io_x_paa(tlb_entries_barrier_9_io_x_paa),
    .io_x_eff(tlb_entries_barrier_9_io_x_eff),
    .io_x_c(tlb_entries_barrier_9_io_x_c),
    .io_y_ppn(tlb_entries_barrier_9_io_y_ppn),
    .io_y_u(tlb_entries_barrier_9_io_y_u),
    .io_y_ae(tlb_entries_barrier_9_io_y_ae),
    .io_y_sw(tlb_entries_barrier_9_io_y_sw),
    .io_y_sx(tlb_entries_barrier_9_io_y_sx),
    .io_y_sr(tlb_entries_barrier_9_io_y_sr),
    .io_y_pw(tlb_entries_barrier_9_io_y_pw),
    .io_y_px(tlb_entries_barrier_9_io_y_px),
    .io_y_pr(tlb_entries_barrier_9_io_y_pr),
    .io_y_ppp(tlb_entries_barrier_9_io_y_ppp),
    .io_y_pal(tlb_entries_barrier_9_io_y_pal),
    .io_y_paa(tlb_entries_barrier_9_io_y_paa),
    .io_y_eff(tlb_entries_barrier_9_io_y_eff),
    .io_y_c(tlb_entries_barrier_9_io_y_c)
  );
  OptimizationBarrier tlb_entries_barrier_10 ( // @[package.scala 236:25]
    .io_x_ppn(tlb_entries_barrier_10_io_x_ppn),
    .io_x_u(tlb_entries_barrier_10_io_x_u),
    .io_x_ae(tlb_entries_barrier_10_io_x_ae),
    .io_x_sw(tlb_entries_barrier_10_io_x_sw),
    .io_x_sx(tlb_entries_barrier_10_io_x_sx),
    .io_x_sr(tlb_entries_barrier_10_io_x_sr),
    .io_x_pw(tlb_entries_barrier_10_io_x_pw),
    .io_x_px(tlb_entries_barrier_10_io_x_px),
    .io_x_pr(tlb_entries_barrier_10_io_x_pr),
    .io_x_ppp(tlb_entries_barrier_10_io_x_ppp),
    .io_x_pal(tlb_entries_barrier_10_io_x_pal),
    .io_x_paa(tlb_entries_barrier_10_io_x_paa),
    .io_x_eff(tlb_entries_barrier_10_io_x_eff),
    .io_x_c(tlb_entries_barrier_10_io_x_c),
    .io_y_ppn(tlb_entries_barrier_10_io_y_ppn),
    .io_y_u(tlb_entries_barrier_10_io_y_u),
    .io_y_ae(tlb_entries_barrier_10_io_y_ae),
    .io_y_sw(tlb_entries_barrier_10_io_y_sw),
    .io_y_sx(tlb_entries_barrier_10_io_y_sx),
    .io_y_sr(tlb_entries_barrier_10_io_y_sr),
    .io_y_pw(tlb_entries_barrier_10_io_y_pw),
    .io_y_px(tlb_entries_barrier_10_io_y_px),
    .io_y_pr(tlb_entries_barrier_10_io_y_pr),
    .io_y_ppp(tlb_entries_barrier_10_io_y_ppp),
    .io_y_pal(tlb_entries_barrier_10_io_y_pal),
    .io_y_paa(tlb_entries_barrier_10_io_y_paa),
    .io_y_eff(tlb_entries_barrier_10_io_y_eff),
    .io_y_c(tlb_entries_barrier_10_io_y_c)
  );
  OptimizationBarrier tlb_entries_barrier_11 ( // @[package.scala 236:25]
    .io_x_ppn(tlb_entries_barrier_11_io_x_ppn),
    .io_x_u(tlb_entries_barrier_11_io_x_u),
    .io_x_ae(tlb_entries_barrier_11_io_x_ae),
    .io_x_sw(tlb_entries_barrier_11_io_x_sw),
    .io_x_sx(tlb_entries_barrier_11_io_x_sx),
    .io_x_sr(tlb_entries_barrier_11_io_x_sr),
    .io_x_pw(tlb_entries_barrier_11_io_x_pw),
    .io_x_px(tlb_entries_barrier_11_io_x_px),
    .io_x_pr(tlb_entries_barrier_11_io_x_pr),
    .io_x_ppp(tlb_entries_barrier_11_io_x_ppp),
    .io_x_pal(tlb_entries_barrier_11_io_x_pal),
    .io_x_paa(tlb_entries_barrier_11_io_x_paa),
    .io_x_eff(tlb_entries_barrier_11_io_x_eff),
    .io_x_c(tlb_entries_barrier_11_io_x_c),
    .io_y_ppn(tlb_entries_barrier_11_io_y_ppn),
    .io_y_u(tlb_entries_barrier_11_io_y_u),
    .io_y_ae(tlb_entries_barrier_11_io_y_ae),
    .io_y_sw(tlb_entries_barrier_11_io_y_sw),
    .io_y_sx(tlb_entries_barrier_11_io_y_sx),
    .io_y_sr(tlb_entries_barrier_11_io_y_sr),
    .io_y_pw(tlb_entries_barrier_11_io_y_pw),
    .io_y_px(tlb_entries_barrier_11_io_y_px),
    .io_y_pr(tlb_entries_barrier_11_io_y_pr),
    .io_y_ppp(tlb_entries_barrier_11_io_y_ppp),
    .io_y_pal(tlb_entries_barrier_11_io_y_pal),
    .io_y_paa(tlb_entries_barrier_11_io_y_paa),
    .io_y_eff(tlb_entries_barrier_11_io_y_eff),
    .io_y_c(tlb_entries_barrier_11_io_y_c)
  );
  OptimizationBarrier tlb_entries_barrier_12 ( // @[package.scala 236:25]
    .io_x_ppn(tlb_entries_barrier_12_io_x_ppn),
    .io_x_u(tlb_entries_barrier_12_io_x_u),
    .io_x_ae(tlb_entries_barrier_12_io_x_ae),
    .io_x_sw(tlb_entries_barrier_12_io_x_sw),
    .io_x_sx(tlb_entries_barrier_12_io_x_sx),
    .io_x_sr(tlb_entries_barrier_12_io_x_sr),
    .io_x_pw(tlb_entries_barrier_12_io_x_pw),
    .io_x_px(tlb_entries_barrier_12_io_x_px),
    .io_x_pr(tlb_entries_barrier_12_io_x_pr),
    .io_x_ppp(tlb_entries_barrier_12_io_x_ppp),
    .io_x_pal(tlb_entries_barrier_12_io_x_pal),
    .io_x_paa(tlb_entries_barrier_12_io_x_paa),
    .io_x_eff(tlb_entries_barrier_12_io_x_eff),
    .io_x_c(tlb_entries_barrier_12_io_x_c),
    .io_y_ppn(tlb_entries_barrier_12_io_y_ppn),
    .io_y_u(tlb_entries_barrier_12_io_y_u),
    .io_y_ae(tlb_entries_barrier_12_io_y_ae),
    .io_y_sw(tlb_entries_barrier_12_io_y_sw),
    .io_y_sx(tlb_entries_barrier_12_io_y_sx),
    .io_y_sr(tlb_entries_barrier_12_io_y_sr),
    .io_y_pw(tlb_entries_barrier_12_io_y_pw),
    .io_y_px(tlb_entries_barrier_12_io_y_px),
    .io_y_pr(tlb_entries_barrier_12_io_y_pr),
    .io_y_ppp(tlb_entries_barrier_12_io_y_ppp),
    .io_y_pal(tlb_entries_barrier_12_io_y_pal),
    .io_y_paa(tlb_entries_barrier_12_io_y_paa),
    .io_y_eff(tlb_entries_barrier_12_io_y_eff),
    .io_y_c(tlb_entries_barrier_12_io_y_c)
  );
  OptimizationBarrier tlb_normal_entries_barrier ( // @[package.scala 236:25]
    .io_x_ppn(tlb_normal_entries_barrier_io_x_ppn),
    .io_x_u(tlb_normal_entries_barrier_io_x_u),
    .io_x_ae(tlb_normal_entries_barrier_io_x_ae),
    .io_x_sw(tlb_normal_entries_barrier_io_x_sw),
    .io_x_sx(tlb_normal_entries_barrier_io_x_sx),
    .io_x_sr(tlb_normal_entries_barrier_io_x_sr),
    .io_x_pw(tlb_normal_entries_barrier_io_x_pw),
    .io_x_px(tlb_normal_entries_barrier_io_x_px),
    .io_x_pr(tlb_normal_entries_barrier_io_x_pr),
    .io_x_ppp(tlb_normal_entries_barrier_io_x_ppp),
    .io_x_pal(tlb_normal_entries_barrier_io_x_pal),
    .io_x_paa(tlb_normal_entries_barrier_io_x_paa),
    .io_x_eff(tlb_normal_entries_barrier_io_x_eff),
    .io_x_c(tlb_normal_entries_barrier_io_x_c),
    .io_y_ppn(tlb_normal_entries_barrier_io_y_ppn),
    .io_y_u(tlb_normal_entries_barrier_io_y_u),
    .io_y_ae(tlb_normal_entries_barrier_io_y_ae),
    .io_y_sw(tlb_normal_entries_barrier_io_y_sw),
    .io_y_sx(tlb_normal_entries_barrier_io_y_sx),
    .io_y_sr(tlb_normal_entries_barrier_io_y_sr),
    .io_y_pw(tlb_normal_entries_barrier_io_y_pw),
    .io_y_px(tlb_normal_entries_barrier_io_y_px),
    .io_y_pr(tlb_normal_entries_barrier_io_y_pr),
    .io_y_ppp(tlb_normal_entries_barrier_io_y_ppp),
    .io_y_pal(tlb_normal_entries_barrier_io_y_pal),
    .io_y_paa(tlb_normal_entries_barrier_io_y_paa),
    .io_y_eff(tlb_normal_entries_barrier_io_y_eff),
    .io_y_c(tlb_normal_entries_barrier_io_y_c)
  );
  OptimizationBarrier tlb_normal_entries_barrier_1 ( // @[package.scala 236:25]
    .io_x_ppn(tlb_normal_entries_barrier_1_io_x_ppn),
    .io_x_u(tlb_normal_entries_barrier_1_io_x_u),
    .io_x_ae(tlb_normal_entries_barrier_1_io_x_ae),
    .io_x_sw(tlb_normal_entries_barrier_1_io_x_sw),
    .io_x_sx(tlb_normal_entries_barrier_1_io_x_sx),
    .io_x_sr(tlb_normal_entries_barrier_1_io_x_sr),
    .io_x_pw(tlb_normal_entries_barrier_1_io_x_pw),
    .io_x_px(tlb_normal_entries_barrier_1_io_x_px),
    .io_x_pr(tlb_normal_entries_barrier_1_io_x_pr),
    .io_x_ppp(tlb_normal_entries_barrier_1_io_x_ppp),
    .io_x_pal(tlb_normal_entries_barrier_1_io_x_pal),
    .io_x_paa(tlb_normal_entries_barrier_1_io_x_paa),
    .io_x_eff(tlb_normal_entries_barrier_1_io_x_eff),
    .io_x_c(tlb_normal_entries_barrier_1_io_x_c),
    .io_y_ppn(tlb_normal_entries_barrier_1_io_y_ppn),
    .io_y_u(tlb_normal_entries_barrier_1_io_y_u),
    .io_y_ae(tlb_normal_entries_barrier_1_io_y_ae),
    .io_y_sw(tlb_normal_entries_barrier_1_io_y_sw),
    .io_y_sx(tlb_normal_entries_barrier_1_io_y_sx),
    .io_y_sr(tlb_normal_entries_barrier_1_io_y_sr),
    .io_y_pw(tlb_normal_entries_barrier_1_io_y_pw),
    .io_y_px(tlb_normal_entries_barrier_1_io_y_px),
    .io_y_pr(tlb_normal_entries_barrier_1_io_y_pr),
    .io_y_ppp(tlb_normal_entries_barrier_1_io_y_ppp),
    .io_y_pal(tlb_normal_entries_barrier_1_io_y_pal),
    .io_y_paa(tlb_normal_entries_barrier_1_io_y_paa),
    .io_y_eff(tlb_normal_entries_barrier_1_io_y_eff),
    .io_y_c(tlb_normal_entries_barrier_1_io_y_c)
  );
  OptimizationBarrier tlb_normal_entries_barrier_2 ( // @[package.scala 236:25]
    .io_x_ppn(tlb_normal_entries_barrier_2_io_x_ppn),
    .io_x_u(tlb_normal_entries_barrier_2_io_x_u),
    .io_x_ae(tlb_normal_entries_barrier_2_io_x_ae),
    .io_x_sw(tlb_normal_entries_barrier_2_io_x_sw),
    .io_x_sx(tlb_normal_entries_barrier_2_io_x_sx),
    .io_x_sr(tlb_normal_entries_barrier_2_io_x_sr),
    .io_x_pw(tlb_normal_entries_barrier_2_io_x_pw),
    .io_x_px(tlb_normal_entries_barrier_2_io_x_px),
    .io_x_pr(tlb_normal_entries_barrier_2_io_x_pr),
    .io_x_ppp(tlb_normal_entries_barrier_2_io_x_ppp),
    .io_x_pal(tlb_normal_entries_barrier_2_io_x_pal),
    .io_x_paa(tlb_normal_entries_barrier_2_io_x_paa),
    .io_x_eff(tlb_normal_entries_barrier_2_io_x_eff),
    .io_x_c(tlb_normal_entries_barrier_2_io_x_c),
    .io_y_ppn(tlb_normal_entries_barrier_2_io_y_ppn),
    .io_y_u(tlb_normal_entries_barrier_2_io_y_u),
    .io_y_ae(tlb_normal_entries_barrier_2_io_y_ae),
    .io_y_sw(tlb_normal_entries_barrier_2_io_y_sw),
    .io_y_sx(tlb_normal_entries_barrier_2_io_y_sx),
    .io_y_sr(tlb_normal_entries_barrier_2_io_y_sr),
    .io_y_pw(tlb_normal_entries_barrier_2_io_y_pw),
    .io_y_px(tlb_normal_entries_barrier_2_io_y_px),
    .io_y_pr(tlb_normal_entries_barrier_2_io_y_pr),
    .io_y_ppp(tlb_normal_entries_barrier_2_io_y_ppp),
    .io_y_pal(tlb_normal_entries_barrier_2_io_y_pal),
    .io_y_paa(tlb_normal_entries_barrier_2_io_y_paa),
    .io_y_eff(tlb_normal_entries_barrier_2_io_y_eff),
    .io_y_c(tlb_normal_entries_barrier_2_io_y_c)
  );
  OptimizationBarrier tlb_normal_entries_barrier_3 ( // @[package.scala 236:25]
    .io_x_ppn(tlb_normal_entries_barrier_3_io_x_ppn),
    .io_x_u(tlb_normal_entries_barrier_3_io_x_u),
    .io_x_ae(tlb_normal_entries_barrier_3_io_x_ae),
    .io_x_sw(tlb_normal_entries_barrier_3_io_x_sw),
    .io_x_sx(tlb_normal_entries_barrier_3_io_x_sx),
    .io_x_sr(tlb_normal_entries_barrier_3_io_x_sr),
    .io_x_pw(tlb_normal_entries_barrier_3_io_x_pw),
    .io_x_px(tlb_normal_entries_barrier_3_io_x_px),
    .io_x_pr(tlb_normal_entries_barrier_3_io_x_pr),
    .io_x_ppp(tlb_normal_entries_barrier_3_io_x_ppp),
    .io_x_pal(tlb_normal_entries_barrier_3_io_x_pal),
    .io_x_paa(tlb_normal_entries_barrier_3_io_x_paa),
    .io_x_eff(tlb_normal_entries_barrier_3_io_x_eff),
    .io_x_c(tlb_normal_entries_barrier_3_io_x_c),
    .io_y_ppn(tlb_normal_entries_barrier_3_io_y_ppn),
    .io_y_u(tlb_normal_entries_barrier_3_io_y_u),
    .io_y_ae(tlb_normal_entries_barrier_3_io_y_ae),
    .io_y_sw(tlb_normal_entries_barrier_3_io_y_sw),
    .io_y_sx(tlb_normal_entries_barrier_3_io_y_sx),
    .io_y_sr(tlb_normal_entries_barrier_3_io_y_sr),
    .io_y_pw(tlb_normal_entries_barrier_3_io_y_pw),
    .io_y_px(tlb_normal_entries_barrier_3_io_y_px),
    .io_y_pr(tlb_normal_entries_barrier_3_io_y_pr),
    .io_y_ppp(tlb_normal_entries_barrier_3_io_y_ppp),
    .io_y_pal(tlb_normal_entries_barrier_3_io_y_pal),
    .io_y_paa(tlb_normal_entries_barrier_3_io_y_paa),
    .io_y_eff(tlb_normal_entries_barrier_3_io_y_eff),
    .io_y_c(tlb_normal_entries_barrier_3_io_y_c)
  );
  OptimizationBarrier tlb_normal_entries_barrier_4 ( // @[package.scala 236:25]
    .io_x_ppn(tlb_normal_entries_barrier_4_io_x_ppn),
    .io_x_u(tlb_normal_entries_barrier_4_io_x_u),
    .io_x_ae(tlb_normal_entries_barrier_4_io_x_ae),
    .io_x_sw(tlb_normal_entries_barrier_4_io_x_sw),
    .io_x_sx(tlb_normal_entries_barrier_4_io_x_sx),
    .io_x_sr(tlb_normal_entries_barrier_4_io_x_sr),
    .io_x_pw(tlb_normal_entries_barrier_4_io_x_pw),
    .io_x_px(tlb_normal_entries_barrier_4_io_x_px),
    .io_x_pr(tlb_normal_entries_barrier_4_io_x_pr),
    .io_x_ppp(tlb_normal_entries_barrier_4_io_x_ppp),
    .io_x_pal(tlb_normal_entries_barrier_4_io_x_pal),
    .io_x_paa(tlb_normal_entries_barrier_4_io_x_paa),
    .io_x_eff(tlb_normal_entries_barrier_4_io_x_eff),
    .io_x_c(tlb_normal_entries_barrier_4_io_x_c),
    .io_y_ppn(tlb_normal_entries_barrier_4_io_y_ppn),
    .io_y_u(tlb_normal_entries_barrier_4_io_y_u),
    .io_y_ae(tlb_normal_entries_barrier_4_io_y_ae),
    .io_y_sw(tlb_normal_entries_barrier_4_io_y_sw),
    .io_y_sx(tlb_normal_entries_barrier_4_io_y_sx),
    .io_y_sr(tlb_normal_entries_barrier_4_io_y_sr),
    .io_y_pw(tlb_normal_entries_barrier_4_io_y_pw),
    .io_y_px(tlb_normal_entries_barrier_4_io_y_px),
    .io_y_pr(tlb_normal_entries_barrier_4_io_y_pr),
    .io_y_ppp(tlb_normal_entries_barrier_4_io_y_ppp),
    .io_y_pal(tlb_normal_entries_barrier_4_io_y_pal),
    .io_y_paa(tlb_normal_entries_barrier_4_io_y_paa),
    .io_y_eff(tlb_normal_entries_barrier_4_io_y_eff),
    .io_y_c(tlb_normal_entries_barrier_4_io_y_c)
  );
  OptimizationBarrier tlb_normal_entries_barrier_5 ( // @[package.scala 236:25]
    .io_x_ppn(tlb_normal_entries_barrier_5_io_x_ppn),
    .io_x_u(tlb_normal_entries_barrier_5_io_x_u),
    .io_x_ae(tlb_normal_entries_barrier_5_io_x_ae),
    .io_x_sw(tlb_normal_entries_barrier_5_io_x_sw),
    .io_x_sx(tlb_normal_entries_barrier_5_io_x_sx),
    .io_x_sr(tlb_normal_entries_barrier_5_io_x_sr),
    .io_x_pw(tlb_normal_entries_barrier_5_io_x_pw),
    .io_x_px(tlb_normal_entries_barrier_5_io_x_px),
    .io_x_pr(tlb_normal_entries_barrier_5_io_x_pr),
    .io_x_ppp(tlb_normal_entries_barrier_5_io_x_ppp),
    .io_x_pal(tlb_normal_entries_barrier_5_io_x_pal),
    .io_x_paa(tlb_normal_entries_barrier_5_io_x_paa),
    .io_x_eff(tlb_normal_entries_barrier_5_io_x_eff),
    .io_x_c(tlb_normal_entries_barrier_5_io_x_c),
    .io_y_ppn(tlb_normal_entries_barrier_5_io_y_ppn),
    .io_y_u(tlb_normal_entries_barrier_5_io_y_u),
    .io_y_ae(tlb_normal_entries_barrier_5_io_y_ae),
    .io_y_sw(tlb_normal_entries_barrier_5_io_y_sw),
    .io_y_sx(tlb_normal_entries_barrier_5_io_y_sx),
    .io_y_sr(tlb_normal_entries_barrier_5_io_y_sr),
    .io_y_pw(tlb_normal_entries_barrier_5_io_y_pw),
    .io_y_px(tlb_normal_entries_barrier_5_io_y_px),
    .io_y_pr(tlb_normal_entries_barrier_5_io_y_pr),
    .io_y_ppp(tlb_normal_entries_barrier_5_io_y_ppp),
    .io_y_pal(tlb_normal_entries_barrier_5_io_y_pal),
    .io_y_paa(tlb_normal_entries_barrier_5_io_y_paa),
    .io_y_eff(tlb_normal_entries_barrier_5_io_y_eff),
    .io_y_c(tlb_normal_entries_barrier_5_io_y_c)
  );
  OptimizationBarrier tlb_normal_entries_barrier_6 ( // @[package.scala 236:25]
    .io_x_ppn(tlb_normal_entries_barrier_6_io_x_ppn),
    .io_x_u(tlb_normal_entries_barrier_6_io_x_u),
    .io_x_ae(tlb_normal_entries_barrier_6_io_x_ae),
    .io_x_sw(tlb_normal_entries_barrier_6_io_x_sw),
    .io_x_sx(tlb_normal_entries_barrier_6_io_x_sx),
    .io_x_sr(tlb_normal_entries_barrier_6_io_x_sr),
    .io_x_pw(tlb_normal_entries_barrier_6_io_x_pw),
    .io_x_px(tlb_normal_entries_barrier_6_io_x_px),
    .io_x_pr(tlb_normal_entries_barrier_6_io_x_pr),
    .io_x_ppp(tlb_normal_entries_barrier_6_io_x_ppp),
    .io_x_pal(tlb_normal_entries_barrier_6_io_x_pal),
    .io_x_paa(tlb_normal_entries_barrier_6_io_x_paa),
    .io_x_eff(tlb_normal_entries_barrier_6_io_x_eff),
    .io_x_c(tlb_normal_entries_barrier_6_io_x_c),
    .io_y_ppn(tlb_normal_entries_barrier_6_io_y_ppn),
    .io_y_u(tlb_normal_entries_barrier_6_io_y_u),
    .io_y_ae(tlb_normal_entries_barrier_6_io_y_ae),
    .io_y_sw(tlb_normal_entries_barrier_6_io_y_sw),
    .io_y_sx(tlb_normal_entries_barrier_6_io_y_sx),
    .io_y_sr(tlb_normal_entries_barrier_6_io_y_sr),
    .io_y_pw(tlb_normal_entries_barrier_6_io_y_pw),
    .io_y_px(tlb_normal_entries_barrier_6_io_y_px),
    .io_y_pr(tlb_normal_entries_barrier_6_io_y_pr),
    .io_y_ppp(tlb_normal_entries_barrier_6_io_y_ppp),
    .io_y_pal(tlb_normal_entries_barrier_6_io_y_pal),
    .io_y_paa(tlb_normal_entries_barrier_6_io_y_paa),
    .io_y_eff(tlb_normal_entries_barrier_6_io_y_eff),
    .io_y_c(tlb_normal_entries_barrier_6_io_y_c)
  );
  OptimizationBarrier tlb_normal_entries_barrier_7 ( // @[package.scala 236:25]
    .io_x_ppn(tlb_normal_entries_barrier_7_io_x_ppn),
    .io_x_u(tlb_normal_entries_barrier_7_io_x_u),
    .io_x_ae(tlb_normal_entries_barrier_7_io_x_ae),
    .io_x_sw(tlb_normal_entries_barrier_7_io_x_sw),
    .io_x_sx(tlb_normal_entries_barrier_7_io_x_sx),
    .io_x_sr(tlb_normal_entries_barrier_7_io_x_sr),
    .io_x_pw(tlb_normal_entries_barrier_7_io_x_pw),
    .io_x_px(tlb_normal_entries_barrier_7_io_x_px),
    .io_x_pr(tlb_normal_entries_barrier_7_io_x_pr),
    .io_x_ppp(tlb_normal_entries_barrier_7_io_x_ppp),
    .io_x_pal(tlb_normal_entries_barrier_7_io_x_pal),
    .io_x_paa(tlb_normal_entries_barrier_7_io_x_paa),
    .io_x_eff(tlb_normal_entries_barrier_7_io_x_eff),
    .io_x_c(tlb_normal_entries_barrier_7_io_x_c),
    .io_y_ppn(tlb_normal_entries_barrier_7_io_y_ppn),
    .io_y_u(tlb_normal_entries_barrier_7_io_y_u),
    .io_y_ae(tlb_normal_entries_barrier_7_io_y_ae),
    .io_y_sw(tlb_normal_entries_barrier_7_io_y_sw),
    .io_y_sx(tlb_normal_entries_barrier_7_io_y_sx),
    .io_y_sr(tlb_normal_entries_barrier_7_io_y_sr),
    .io_y_pw(tlb_normal_entries_barrier_7_io_y_pw),
    .io_y_px(tlb_normal_entries_barrier_7_io_y_px),
    .io_y_pr(tlb_normal_entries_barrier_7_io_y_pr),
    .io_y_ppp(tlb_normal_entries_barrier_7_io_y_ppp),
    .io_y_pal(tlb_normal_entries_barrier_7_io_y_pal),
    .io_y_paa(tlb_normal_entries_barrier_7_io_y_paa),
    .io_y_eff(tlb_normal_entries_barrier_7_io_y_eff),
    .io_y_c(tlb_normal_entries_barrier_7_io_y_c)
  );
  OptimizationBarrier tlb_normal_entries_barrier_8 ( // @[package.scala 236:25]
    .io_x_ppn(tlb_normal_entries_barrier_8_io_x_ppn),
    .io_x_u(tlb_normal_entries_barrier_8_io_x_u),
    .io_x_ae(tlb_normal_entries_barrier_8_io_x_ae),
    .io_x_sw(tlb_normal_entries_barrier_8_io_x_sw),
    .io_x_sx(tlb_normal_entries_barrier_8_io_x_sx),
    .io_x_sr(tlb_normal_entries_barrier_8_io_x_sr),
    .io_x_pw(tlb_normal_entries_barrier_8_io_x_pw),
    .io_x_px(tlb_normal_entries_barrier_8_io_x_px),
    .io_x_pr(tlb_normal_entries_barrier_8_io_x_pr),
    .io_x_ppp(tlb_normal_entries_barrier_8_io_x_ppp),
    .io_x_pal(tlb_normal_entries_barrier_8_io_x_pal),
    .io_x_paa(tlb_normal_entries_barrier_8_io_x_paa),
    .io_x_eff(tlb_normal_entries_barrier_8_io_x_eff),
    .io_x_c(tlb_normal_entries_barrier_8_io_x_c),
    .io_y_ppn(tlb_normal_entries_barrier_8_io_y_ppn),
    .io_y_u(tlb_normal_entries_barrier_8_io_y_u),
    .io_y_ae(tlb_normal_entries_barrier_8_io_y_ae),
    .io_y_sw(tlb_normal_entries_barrier_8_io_y_sw),
    .io_y_sx(tlb_normal_entries_barrier_8_io_y_sx),
    .io_y_sr(tlb_normal_entries_barrier_8_io_y_sr),
    .io_y_pw(tlb_normal_entries_barrier_8_io_y_pw),
    .io_y_px(tlb_normal_entries_barrier_8_io_y_px),
    .io_y_pr(tlb_normal_entries_barrier_8_io_y_pr),
    .io_y_ppp(tlb_normal_entries_barrier_8_io_y_ppp),
    .io_y_pal(tlb_normal_entries_barrier_8_io_y_pal),
    .io_y_paa(tlb_normal_entries_barrier_8_io_y_paa),
    .io_y_eff(tlb_normal_entries_barrier_8_io_y_eff),
    .io_y_c(tlb_normal_entries_barrier_8_io_y_c)
  );
  OptimizationBarrier tlb_normal_entries_barrier_9 ( // @[package.scala 236:25]
    .io_x_ppn(tlb_normal_entries_barrier_9_io_x_ppn),
    .io_x_u(tlb_normal_entries_barrier_9_io_x_u),
    .io_x_ae(tlb_normal_entries_barrier_9_io_x_ae),
    .io_x_sw(tlb_normal_entries_barrier_9_io_x_sw),
    .io_x_sx(tlb_normal_entries_barrier_9_io_x_sx),
    .io_x_sr(tlb_normal_entries_barrier_9_io_x_sr),
    .io_x_pw(tlb_normal_entries_barrier_9_io_x_pw),
    .io_x_px(tlb_normal_entries_barrier_9_io_x_px),
    .io_x_pr(tlb_normal_entries_barrier_9_io_x_pr),
    .io_x_ppp(tlb_normal_entries_barrier_9_io_x_ppp),
    .io_x_pal(tlb_normal_entries_barrier_9_io_x_pal),
    .io_x_paa(tlb_normal_entries_barrier_9_io_x_paa),
    .io_x_eff(tlb_normal_entries_barrier_9_io_x_eff),
    .io_x_c(tlb_normal_entries_barrier_9_io_x_c),
    .io_y_ppn(tlb_normal_entries_barrier_9_io_y_ppn),
    .io_y_u(tlb_normal_entries_barrier_9_io_y_u),
    .io_y_ae(tlb_normal_entries_barrier_9_io_y_ae),
    .io_y_sw(tlb_normal_entries_barrier_9_io_y_sw),
    .io_y_sx(tlb_normal_entries_barrier_9_io_y_sx),
    .io_y_sr(tlb_normal_entries_barrier_9_io_y_sr),
    .io_y_pw(tlb_normal_entries_barrier_9_io_y_pw),
    .io_y_px(tlb_normal_entries_barrier_9_io_y_px),
    .io_y_pr(tlb_normal_entries_barrier_9_io_y_pr),
    .io_y_ppp(tlb_normal_entries_barrier_9_io_y_ppp),
    .io_y_pal(tlb_normal_entries_barrier_9_io_y_pal),
    .io_y_paa(tlb_normal_entries_barrier_9_io_y_paa),
    .io_y_eff(tlb_normal_entries_barrier_9_io_y_eff),
    .io_y_c(tlb_normal_entries_barrier_9_io_y_c)
  );
  OptimizationBarrier tlb_normal_entries_barrier_10 ( // @[package.scala 236:25]
    .io_x_ppn(tlb_normal_entries_barrier_10_io_x_ppn),
    .io_x_u(tlb_normal_entries_barrier_10_io_x_u),
    .io_x_ae(tlb_normal_entries_barrier_10_io_x_ae),
    .io_x_sw(tlb_normal_entries_barrier_10_io_x_sw),
    .io_x_sx(tlb_normal_entries_barrier_10_io_x_sx),
    .io_x_sr(tlb_normal_entries_barrier_10_io_x_sr),
    .io_x_pw(tlb_normal_entries_barrier_10_io_x_pw),
    .io_x_px(tlb_normal_entries_barrier_10_io_x_px),
    .io_x_pr(tlb_normal_entries_barrier_10_io_x_pr),
    .io_x_ppp(tlb_normal_entries_barrier_10_io_x_ppp),
    .io_x_pal(tlb_normal_entries_barrier_10_io_x_pal),
    .io_x_paa(tlb_normal_entries_barrier_10_io_x_paa),
    .io_x_eff(tlb_normal_entries_barrier_10_io_x_eff),
    .io_x_c(tlb_normal_entries_barrier_10_io_x_c),
    .io_y_ppn(tlb_normal_entries_barrier_10_io_y_ppn),
    .io_y_u(tlb_normal_entries_barrier_10_io_y_u),
    .io_y_ae(tlb_normal_entries_barrier_10_io_y_ae),
    .io_y_sw(tlb_normal_entries_barrier_10_io_y_sw),
    .io_y_sx(tlb_normal_entries_barrier_10_io_y_sx),
    .io_y_sr(tlb_normal_entries_barrier_10_io_y_sr),
    .io_y_pw(tlb_normal_entries_barrier_10_io_y_pw),
    .io_y_px(tlb_normal_entries_barrier_10_io_y_px),
    .io_y_pr(tlb_normal_entries_barrier_10_io_y_pr),
    .io_y_ppp(tlb_normal_entries_barrier_10_io_y_ppp),
    .io_y_pal(tlb_normal_entries_barrier_10_io_y_pal),
    .io_y_paa(tlb_normal_entries_barrier_10_io_y_paa),
    .io_y_eff(tlb_normal_entries_barrier_10_io_y_eff),
    .io_y_c(tlb_normal_entries_barrier_10_io_y_c)
  );
  OptimizationBarrier tlb_normal_entries_barrier_11 ( // @[package.scala 236:25]
    .io_x_ppn(tlb_normal_entries_barrier_11_io_x_ppn),
    .io_x_u(tlb_normal_entries_barrier_11_io_x_u),
    .io_x_ae(tlb_normal_entries_barrier_11_io_x_ae),
    .io_x_sw(tlb_normal_entries_barrier_11_io_x_sw),
    .io_x_sx(tlb_normal_entries_barrier_11_io_x_sx),
    .io_x_sr(tlb_normal_entries_barrier_11_io_x_sr),
    .io_x_pw(tlb_normal_entries_barrier_11_io_x_pw),
    .io_x_px(tlb_normal_entries_barrier_11_io_x_px),
    .io_x_pr(tlb_normal_entries_barrier_11_io_x_pr),
    .io_x_ppp(tlb_normal_entries_barrier_11_io_x_ppp),
    .io_x_pal(tlb_normal_entries_barrier_11_io_x_pal),
    .io_x_paa(tlb_normal_entries_barrier_11_io_x_paa),
    .io_x_eff(tlb_normal_entries_barrier_11_io_x_eff),
    .io_x_c(tlb_normal_entries_barrier_11_io_x_c),
    .io_y_ppn(tlb_normal_entries_barrier_11_io_y_ppn),
    .io_y_u(tlb_normal_entries_barrier_11_io_y_u),
    .io_y_ae(tlb_normal_entries_barrier_11_io_y_ae),
    .io_y_sw(tlb_normal_entries_barrier_11_io_y_sw),
    .io_y_sx(tlb_normal_entries_barrier_11_io_y_sx),
    .io_y_sr(tlb_normal_entries_barrier_11_io_y_sr),
    .io_y_pw(tlb_normal_entries_barrier_11_io_y_pw),
    .io_y_px(tlb_normal_entries_barrier_11_io_y_px),
    .io_y_pr(tlb_normal_entries_barrier_11_io_y_pr),
    .io_y_ppp(tlb_normal_entries_barrier_11_io_y_ppp),
    .io_y_pal(tlb_normal_entries_barrier_11_io_y_pal),
    .io_y_paa(tlb_normal_entries_barrier_11_io_y_paa),
    .io_y_eff(tlb_normal_entries_barrier_11_io_y_eff),
    .io_y_c(tlb_normal_entries_barrier_11_io_y_c)
  );
  OptimizationBarrier pma_checker_mpu_ppn_data_barrier ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_mpu_ppn_data_barrier_io_x_ppn),
    .io_x_u(pma_checker_mpu_ppn_data_barrier_io_x_u),
    .io_x_ae(pma_checker_mpu_ppn_data_barrier_io_x_ae),
    .io_x_sw(pma_checker_mpu_ppn_data_barrier_io_x_sw),
    .io_x_sx(pma_checker_mpu_ppn_data_barrier_io_x_sx),
    .io_x_sr(pma_checker_mpu_ppn_data_barrier_io_x_sr),
    .io_x_pw(pma_checker_mpu_ppn_data_barrier_io_x_pw),
    .io_x_px(pma_checker_mpu_ppn_data_barrier_io_x_px),
    .io_x_pr(pma_checker_mpu_ppn_data_barrier_io_x_pr),
    .io_x_ppp(pma_checker_mpu_ppn_data_barrier_io_x_ppp),
    .io_x_pal(pma_checker_mpu_ppn_data_barrier_io_x_pal),
    .io_x_paa(pma_checker_mpu_ppn_data_barrier_io_x_paa),
    .io_x_eff(pma_checker_mpu_ppn_data_barrier_io_x_eff),
    .io_x_c(pma_checker_mpu_ppn_data_barrier_io_x_c),
    .io_y_ppn(pma_checker_mpu_ppn_data_barrier_io_y_ppn),
    .io_y_u(pma_checker_mpu_ppn_data_barrier_io_y_u),
    .io_y_ae(pma_checker_mpu_ppn_data_barrier_io_y_ae),
    .io_y_sw(pma_checker_mpu_ppn_data_barrier_io_y_sw),
    .io_y_sx(pma_checker_mpu_ppn_data_barrier_io_y_sx),
    .io_y_sr(pma_checker_mpu_ppn_data_barrier_io_y_sr),
    .io_y_pw(pma_checker_mpu_ppn_data_barrier_io_y_pw),
    .io_y_px(pma_checker_mpu_ppn_data_barrier_io_y_px),
    .io_y_pr(pma_checker_mpu_ppn_data_barrier_io_y_pr),
    .io_y_ppp(pma_checker_mpu_ppn_data_barrier_io_y_ppp),
    .io_y_pal(pma_checker_mpu_ppn_data_barrier_io_y_pal),
    .io_y_paa(pma_checker_mpu_ppn_data_barrier_io_y_paa),
    .io_y_eff(pma_checker_mpu_ppn_data_barrier_io_y_eff),
    .io_y_c(pma_checker_mpu_ppn_data_barrier_io_y_c)
  );
  PMPChecker pma_checker_pmp ( // @[TLB.scala 190:19]
    .io_prv(pma_checker_pmp_io_prv),
    .io_pmp_0_cfg_l(pma_checker_pmp_io_pmp_0_cfg_l),
    .io_pmp_0_cfg_a(pma_checker_pmp_io_pmp_0_cfg_a),
    .io_pmp_0_cfg_x(pma_checker_pmp_io_pmp_0_cfg_x),
    .io_pmp_0_cfg_w(pma_checker_pmp_io_pmp_0_cfg_w),
    .io_pmp_0_cfg_r(pma_checker_pmp_io_pmp_0_cfg_r),
    .io_pmp_0_addr(pma_checker_pmp_io_pmp_0_addr),
    .io_pmp_0_mask(pma_checker_pmp_io_pmp_0_mask),
    .io_pmp_1_cfg_l(pma_checker_pmp_io_pmp_1_cfg_l),
    .io_pmp_1_cfg_a(pma_checker_pmp_io_pmp_1_cfg_a),
    .io_pmp_1_cfg_x(pma_checker_pmp_io_pmp_1_cfg_x),
    .io_pmp_1_cfg_w(pma_checker_pmp_io_pmp_1_cfg_w),
    .io_pmp_1_cfg_r(pma_checker_pmp_io_pmp_1_cfg_r),
    .io_pmp_1_addr(pma_checker_pmp_io_pmp_1_addr),
    .io_pmp_1_mask(pma_checker_pmp_io_pmp_1_mask),
    .io_pmp_2_cfg_l(pma_checker_pmp_io_pmp_2_cfg_l),
    .io_pmp_2_cfg_a(pma_checker_pmp_io_pmp_2_cfg_a),
    .io_pmp_2_cfg_x(pma_checker_pmp_io_pmp_2_cfg_x),
    .io_pmp_2_cfg_w(pma_checker_pmp_io_pmp_2_cfg_w),
    .io_pmp_2_cfg_r(pma_checker_pmp_io_pmp_2_cfg_r),
    .io_pmp_2_addr(pma_checker_pmp_io_pmp_2_addr),
    .io_pmp_2_mask(pma_checker_pmp_io_pmp_2_mask),
    .io_pmp_3_cfg_l(pma_checker_pmp_io_pmp_3_cfg_l),
    .io_pmp_3_cfg_a(pma_checker_pmp_io_pmp_3_cfg_a),
    .io_pmp_3_cfg_x(pma_checker_pmp_io_pmp_3_cfg_x),
    .io_pmp_3_cfg_w(pma_checker_pmp_io_pmp_3_cfg_w),
    .io_pmp_3_cfg_r(pma_checker_pmp_io_pmp_3_cfg_r),
    .io_pmp_3_addr(pma_checker_pmp_io_pmp_3_addr),
    .io_pmp_3_mask(pma_checker_pmp_io_pmp_3_mask),
    .io_pmp_4_cfg_l(pma_checker_pmp_io_pmp_4_cfg_l),
    .io_pmp_4_cfg_a(pma_checker_pmp_io_pmp_4_cfg_a),
    .io_pmp_4_cfg_x(pma_checker_pmp_io_pmp_4_cfg_x),
    .io_pmp_4_cfg_w(pma_checker_pmp_io_pmp_4_cfg_w),
    .io_pmp_4_cfg_r(pma_checker_pmp_io_pmp_4_cfg_r),
    .io_pmp_4_addr(pma_checker_pmp_io_pmp_4_addr),
    .io_pmp_4_mask(pma_checker_pmp_io_pmp_4_mask),
    .io_pmp_5_cfg_l(pma_checker_pmp_io_pmp_5_cfg_l),
    .io_pmp_5_cfg_a(pma_checker_pmp_io_pmp_5_cfg_a),
    .io_pmp_5_cfg_x(pma_checker_pmp_io_pmp_5_cfg_x),
    .io_pmp_5_cfg_w(pma_checker_pmp_io_pmp_5_cfg_w),
    .io_pmp_5_cfg_r(pma_checker_pmp_io_pmp_5_cfg_r),
    .io_pmp_5_addr(pma_checker_pmp_io_pmp_5_addr),
    .io_pmp_5_mask(pma_checker_pmp_io_pmp_5_mask),
    .io_pmp_6_cfg_l(pma_checker_pmp_io_pmp_6_cfg_l),
    .io_pmp_6_cfg_a(pma_checker_pmp_io_pmp_6_cfg_a),
    .io_pmp_6_cfg_x(pma_checker_pmp_io_pmp_6_cfg_x),
    .io_pmp_6_cfg_w(pma_checker_pmp_io_pmp_6_cfg_w),
    .io_pmp_6_cfg_r(pma_checker_pmp_io_pmp_6_cfg_r),
    .io_pmp_6_addr(pma_checker_pmp_io_pmp_6_addr),
    .io_pmp_6_mask(pma_checker_pmp_io_pmp_6_mask),
    .io_pmp_7_cfg_l(pma_checker_pmp_io_pmp_7_cfg_l),
    .io_pmp_7_cfg_a(pma_checker_pmp_io_pmp_7_cfg_a),
    .io_pmp_7_cfg_x(pma_checker_pmp_io_pmp_7_cfg_x),
    .io_pmp_7_cfg_w(pma_checker_pmp_io_pmp_7_cfg_w),
    .io_pmp_7_cfg_r(pma_checker_pmp_io_pmp_7_cfg_r),
    .io_pmp_7_addr(pma_checker_pmp_io_pmp_7_addr),
    .io_pmp_7_mask(pma_checker_pmp_io_pmp_7_mask),
    .io_addr(pma_checker_pmp_io_addr),
    .io_size(pma_checker_pmp_io_size),
    .io_r(pma_checker_pmp_io_r),
    .io_w(pma_checker_pmp_io_w),
    .io_x(pma_checker_pmp_io_x)
  );
  OptimizationBarrier pma_checker_ppn_data_barrier ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_ppn_data_barrier_io_x_ppn),
    .io_x_u(pma_checker_ppn_data_barrier_io_x_u),
    .io_x_ae(pma_checker_ppn_data_barrier_io_x_ae),
    .io_x_sw(pma_checker_ppn_data_barrier_io_x_sw),
    .io_x_sx(pma_checker_ppn_data_barrier_io_x_sx),
    .io_x_sr(pma_checker_ppn_data_barrier_io_x_sr),
    .io_x_pw(pma_checker_ppn_data_barrier_io_x_pw),
    .io_x_px(pma_checker_ppn_data_barrier_io_x_px),
    .io_x_pr(pma_checker_ppn_data_barrier_io_x_pr),
    .io_x_ppp(pma_checker_ppn_data_barrier_io_x_ppp),
    .io_x_pal(pma_checker_ppn_data_barrier_io_x_pal),
    .io_x_paa(pma_checker_ppn_data_barrier_io_x_paa),
    .io_x_eff(pma_checker_ppn_data_barrier_io_x_eff),
    .io_x_c(pma_checker_ppn_data_barrier_io_x_c),
    .io_y_ppn(pma_checker_ppn_data_barrier_io_y_ppn),
    .io_y_u(pma_checker_ppn_data_barrier_io_y_u),
    .io_y_ae(pma_checker_ppn_data_barrier_io_y_ae),
    .io_y_sw(pma_checker_ppn_data_barrier_io_y_sw),
    .io_y_sx(pma_checker_ppn_data_barrier_io_y_sx),
    .io_y_sr(pma_checker_ppn_data_barrier_io_y_sr),
    .io_y_pw(pma_checker_ppn_data_barrier_io_y_pw),
    .io_y_px(pma_checker_ppn_data_barrier_io_y_px),
    .io_y_pr(pma_checker_ppn_data_barrier_io_y_pr),
    .io_y_ppp(pma_checker_ppn_data_barrier_io_y_ppp),
    .io_y_pal(pma_checker_ppn_data_barrier_io_y_pal),
    .io_y_paa(pma_checker_ppn_data_barrier_io_y_paa),
    .io_y_eff(pma_checker_ppn_data_barrier_io_y_eff),
    .io_y_c(pma_checker_ppn_data_barrier_io_y_c)
  );
  OptimizationBarrier pma_checker_ppn_data_barrier_1 ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_ppn_data_barrier_1_io_x_ppn),
    .io_x_u(pma_checker_ppn_data_barrier_1_io_x_u),
    .io_x_ae(pma_checker_ppn_data_barrier_1_io_x_ae),
    .io_x_sw(pma_checker_ppn_data_barrier_1_io_x_sw),
    .io_x_sx(pma_checker_ppn_data_barrier_1_io_x_sx),
    .io_x_sr(pma_checker_ppn_data_barrier_1_io_x_sr),
    .io_x_pw(pma_checker_ppn_data_barrier_1_io_x_pw),
    .io_x_px(pma_checker_ppn_data_barrier_1_io_x_px),
    .io_x_pr(pma_checker_ppn_data_barrier_1_io_x_pr),
    .io_x_ppp(pma_checker_ppn_data_barrier_1_io_x_ppp),
    .io_x_pal(pma_checker_ppn_data_barrier_1_io_x_pal),
    .io_x_paa(pma_checker_ppn_data_barrier_1_io_x_paa),
    .io_x_eff(pma_checker_ppn_data_barrier_1_io_x_eff),
    .io_x_c(pma_checker_ppn_data_barrier_1_io_x_c),
    .io_y_ppn(pma_checker_ppn_data_barrier_1_io_y_ppn),
    .io_y_u(pma_checker_ppn_data_barrier_1_io_y_u),
    .io_y_ae(pma_checker_ppn_data_barrier_1_io_y_ae),
    .io_y_sw(pma_checker_ppn_data_barrier_1_io_y_sw),
    .io_y_sx(pma_checker_ppn_data_barrier_1_io_y_sx),
    .io_y_sr(pma_checker_ppn_data_barrier_1_io_y_sr),
    .io_y_pw(pma_checker_ppn_data_barrier_1_io_y_pw),
    .io_y_px(pma_checker_ppn_data_barrier_1_io_y_px),
    .io_y_pr(pma_checker_ppn_data_barrier_1_io_y_pr),
    .io_y_ppp(pma_checker_ppn_data_barrier_1_io_y_ppp),
    .io_y_pal(pma_checker_ppn_data_barrier_1_io_y_pal),
    .io_y_paa(pma_checker_ppn_data_barrier_1_io_y_paa),
    .io_y_eff(pma_checker_ppn_data_barrier_1_io_y_eff),
    .io_y_c(pma_checker_ppn_data_barrier_1_io_y_c)
  );
  OptimizationBarrier pma_checker_ppn_data_barrier_2 ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_ppn_data_barrier_2_io_x_ppn),
    .io_x_u(pma_checker_ppn_data_barrier_2_io_x_u),
    .io_x_ae(pma_checker_ppn_data_barrier_2_io_x_ae),
    .io_x_sw(pma_checker_ppn_data_barrier_2_io_x_sw),
    .io_x_sx(pma_checker_ppn_data_barrier_2_io_x_sx),
    .io_x_sr(pma_checker_ppn_data_barrier_2_io_x_sr),
    .io_x_pw(pma_checker_ppn_data_barrier_2_io_x_pw),
    .io_x_px(pma_checker_ppn_data_barrier_2_io_x_px),
    .io_x_pr(pma_checker_ppn_data_barrier_2_io_x_pr),
    .io_x_ppp(pma_checker_ppn_data_barrier_2_io_x_ppp),
    .io_x_pal(pma_checker_ppn_data_barrier_2_io_x_pal),
    .io_x_paa(pma_checker_ppn_data_barrier_2_io_x_paa),
    .io_x_eff(pma_checker_ppn_data_barrier_2_io_x_eff),
    .io_x_c(pma_checker_ppn_data_barrier_2_io_x_c),
    .io_y_ppn(pma_checker_ppn_data_barrier_2_io_y_ppn),
    .io_y_u(pma_checker_ppn_data_barrier_2_io_y_u),
    .io_y_ae(pma_checker_ppn_data_barrier_2_io_y_ae),
    .io_y_sw(pma_checker_ppn_data_barrier_2_io_y_sw),
    .io_y_sx(pma_checker_ppn_data_barrier_2_io_y_sx),
    .io_y_sr(pma_checker_ppn_data_barrier_2_io_y_sr),
    .io_y_pw(pma_checker_ppn_data_barrier_2_io_y_pw),
    .io_y_px(pma_checker_ppn_data_barrier_2_io_y_px),
    .io_y_pr(pma_checker_ppn_data_barrier_2_io_y_pr),
    .io_y_ppp(pma_checker_ppn_data_barrier_2_io_y_ppp),
    .io_y_pal(pma_checker_ppn_data_barrier_2_io_y_pal),
    .io_y_paa(pma_checker_ppn_data_barrier_2_io_y_paa),
    .io_y_eff(pma_checker_ppn_data_barrier_2_io_y_eff),
    .io_y_c(pma_checker_ppn_data_barrier_2_io_y_c)
  );
  OptimizationBarrier pma_checker_ppn_data_barrier_3 ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_ppn_data_barrier_3_io_x_ppn),
    .io_x_u(pma_checker_ppn_data_barrier_3_io_x_u),
    .io_x_ae(pma_checker_ppn_data_barrier_3_io_x_ae),
    .io_x_sw(pma_checker_ppn_data_barrier_3_io_x_sw),
    .io_x_sx(pma_checker_ppn_data_barrier_3_io_x_sx),
    .io_x_sr(pma_checker_ppn_data_barrier_3_io_x_sr),
    .io_x_pw(pma_checker_ppn_data_barrier_3_io_x_pw),
    .io_x_px(pma_checker_ppn_data_barrier_3_io_x_px),
    .io_x_pr(pma_checker_ppn_data_barrier_3_io_x_pr),
    .io_x_ppp(pma_checker_ppn_data_barrier_3_io_x_ppp),
    .io_x_pal(pma_checker_ppn_data_barrier_3_io_x_pal),
    .io_x_paa(pma_checker_ppn_data_barrier_3_io_x_paa),
    .io_x_eff(pma_checker_ppn_data_barrier_3_io_x_eff),
    .io_x_c(pma_checker_ppn_data_barrier_3_io_x_c),
    .io_y_ppn(pma_checker_ppn_data_barrier_3_io_y_ppn),
    .io_y_u(pma_checker_ppn_data_barrier_3_io_y_u),
    .io_y_ae(pma_checker_ppn_data_barrier_3_io_y_ae),
    .io_y_sw(pma_checker_ppn_data_barrier_3_io_y_sw),
    .io_y_sx(pma_checker_ppn_data_barrier_3_io_y_sx),
    .io_y_sr(pma_checker_ppn_data_barrier_3_io_y_sr),
    .io_y_pw(pma_checker_ppn_data_barrier_3_io_y_pw),
    .io_y_px(pma_checker_ppn_data_barrier_3_io_y_px),
    .io_y_pr(pma_checker_ppn_data_barrier_3_io_y_pr),
    .io_y_ppp(pma_checker_ppn_data_barrier_3_io_y_ppp),
    .io_y_pal(pma_checker_ppn_data_barrier_3_io_y_pal),
    .io_y_paa(pma_checker_ppn_data_barrier_3_io_y_paa),
    .io_y_eff(pma_checker_ppn_data_barrier_3_io_y_eff),
    .io_y_c(pma_checker_ppn_data_barrier_3_io_y_c)
  );
  OptimizationBarrier pma_checker_ppn_data_barrier_4 ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_ppn_data_barrier_4_io_x_ppn),
    .io_x_u(pma_checker_ppn_data_barrier_4_io_x_u),
    .io_x_ae(pma_checker_ppn_data_barrier_4_io_x_ae),
    .io_x_sw(pma_checker_ppn_data_barrier_4_io_x_sw),
    .io_x_sx(pma_checker_ppn_data_barrier_4_io_x_sx),
    .io_x_sr(pma_checker_ppn_data_barrier_4_io_x_sr),
    .io_x_pw(pma_checker_ppn_data_barrier_4_io_x_pw),
    .io_x_px(pma_checker_ppn_data_barrier_4_io_x_px),
    .io_x_pr(pma_checker_ppn_data_barrier_4_io_x_pr),
    .io_x_ppp(pma_checker_ppn_data_barrier_4_io_x_ppp),
    .io_x_pal(pma_checker_ppn_data_barrier_4_io_x_pal),
    .io_x_paa(pma_checker_ppn_data_barrier_4_io_x_paa),
    .io_x_eff(pma_checker_ppn_data_barrier_4_io_x_eff),
    .io_x_c(pma_checker_ppn_data_barrier_4_io_x_c),
    .io_y_ppn(pma_checker_ppn_data_barrier_4_io_y_ppn),
    .io_y_u(pma_checker_ppn_data_barrier_4_io_y_u),
    .io_y_ae(pma_checker_ppn_data_barrier_4_io_y_ae),
    .io_y_sw(pma_checker_ppn_data_barrier_4_io_y_sw),
    .io_y_sx(pma_checker_ppn_data_barrier_4_io_y_sx),
    .io_y_sr(pma_checker_ppn_data_barrier_4_io_y_sr),
    .io_y_pw(pma_checker_ppn_data_barrier_4_io_y_pw),
    .io_y_px(pma_checker_ppn_data_barrier_4_io_y_px),
    .io_y_pr(pma_checker_ppn_data_barrier_4_io_y_pr),
    .io_y_ppp(pma_checker_ppn_data_barrier_4_io_y_ppp),
    .io_y_pal(pma_checker_ppn_data_barrier_4_io_y_pal),
    .io_y_paa(pma_checker_ppn_data_barrier_4_io_y_paa),
    .io_y_eff(pma_checker_ppn_data_barrier_4_io_y_eff),
    .io_y_c(pma_checker_ppn_data_barrier_4_io_y_c)
  );
  OptimizationBarrier pma_checker_ppn_data_barrier_5 ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_ppn_data_barrier_5_io_x_ppn),
    .io_x_u(pma_checker_ppn_data_barrier_5_io_x_u),
    .io_x_ae(pma_checker_ppn_data_barrier_5_io_x_ae),
    .io_x_sw(pma_checker_ppn_data_barrier_5_io_x_sw),
    .io_x_sx(pma_checker_ppn_data_barrier_5_io_x_sx),
    .io_x_sr(pma_checker_ppn_data_barrier_5_io_x_sr),
    .io_x_pw(pma_checker_ppn_data_barrier_5_io_x_pw),
    .io_x_px(pma_checker_ppn_data_barrier_5_io_x_px),
    .io_x_pr(pma_checker_ppn_data_barrier_5_io_x_pr),
    .io_x_ppp(pma_checker_ppn_data_barrier_5_io_x_ppp),
    .io_x_pal(pma_checker_ppn_data_barrier_5_io_x_pal),
    .io_x_paa(pma_checker_ppn_data_barrier_5_io_x_paa),
    .io_x_eff(pma_checker_ppn_data_barrier_5_io_x_eff),
    .io_x_c(pma_checker_ppn_data_barrier_5_io_x_c),
    .io_y_ppn(pma_checker_ppn_data_barrier_5_io_y_ppn),
    .io_y_u(pma_checker_ppn_data_barrier_5_io_y_u),
    .io_y_ae(pma_checker_ppn_data_barrier_5_io_y_ae),
    .io_y_sw(pma_checker_ppn_data_barrier_5_io_y_sw),
    .io_y_sx(pma_checker_ppn_data_barrier_5_io_y_sx),
    .io_y_sr(pma_checker_ppn_data_barrier_5_io_y_sr),
    .io_y_pw(pma_checker_ppn_data_barrier_5_io_y_pw),
    .io_y_px(pma_checker_ppn_data_barrier_5_io_y_px),
    .io_y_pr(pma_checker_ppn_data_barrier_5_io_y_pr),
    .io_y_ppp(pma_checker_ppn_data_barrier_5_io_y_ppp),
    .io_y_pal(pma_checker_ppn_data_barrier_5_io_y_pal),
    .io_y_paa(pma_checker_ppn_data_barrier_5_io_y_paa),
    .io_y_eff(pma_checker_ppn_data_barrier_5_io_y_eff),
    .io_y_c(pma_checker_ppn_data_barrier_5_io_y_c)
  );
  OptimizationBarrier pma_checker_ppn_data_barrier_6 ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_ppn_data_barrier_6_io_x_ppn),
    .io_x_u(pma_checker_ppn_data_barrier_6_io_x_u),
    .io_x_ae(pma_checker_ppn_data_barrier_6_io_x_ae),
    .io_x_sw(pma_checker_ppn_data_barrier_6_io_x_sw),
    .io_x_sx(pma_checker_ppn_data_barrier_6_io_x_sx),
    .io_x_sr(pma_checker_ppn_data_barrier_6_io_x_sr),
    .io_x_pw(pma_checker_ppn_data_barrier_6_io_x_pw),
    .io_x_px(pma_checker_ppn_data_barrier_6_io_x_px),
    .io_x_pr(pma_checker_ppn_data_barrier_6_io_x_pr),
    .io_x_ppp(pma_checker_ppn_data_barrier_6_io_x_ppp),
    .io_x_pal(pma_checker_ppn_data_barrier_6_io_x_pal),
    .io_x_paa(pma_checker_ppn_data_barrier_6_io_x_paa),
    .io_x_eff(pma_checker_ppn_data_barrier_6_io_x_eff),
    .io_x_c(pma_checker_ppn_data_barrier_6_io_x_c),
    .io_y_ppn(pma_checker_ppn_data_barrier_6_io_y_ppn),
    .io_y_u(pma_checker_ppn_data_barrier_6_io_y_u),
    .io_y_ae(pma_checker_ppn_data_barrier_6_io_y_ae),
    .io_y_sw(pma_checker_ppn_data_barrier_6_io_y_sw),
    .io_y_sx(pma_checker_ppn_data_barrier_6_io_y_sx),
    .io_y_sr(pma_checker_ppn_data_barrier_6_io_y_sr),
    .io_y_pw(pma_checker_ppn_data_barrier_6_io_y_pw),
    .io_y_px(pma_checker_ppn_data_barrier_6_io_y_px),
    .io_y_pr(pma_checker_ppn_data_barrier_6_io_y_pr),
    .io_y_ppp(pma_checker_ppn_data_barrier_6_io_y_ppp),
    .io_y_pal(pma_checker_ppn_data_barrier_6_io_y_pal),
    .io_y_paa(pma_checker_ppn_data_barrier_6_io_y_paa),
    .io_y_eff(pma_checker_ppn_data_barrier_6_io_y_eff),
    .io_y_c(pma_checker_ppn_data_barrier_6_io_y_c)
  );
  OptimizationBarrier pma_checker_ppn_data_barrier_7 ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_ppn_data_barrier_7_io_x_ppn),
    .io_x_u(pma_checker_ppn_data_barrier_7_io_x_u),
    .io_x_ae(pma_checker_ppn_data_barrier_7_io_x_ae),
    .io_x_sw(pma_checker_ppn_data_barrier_7_io_x_sw),
    .io_x_sx(pma_checker_ppn_data_barrier_7_io_x_sx),
    .io_x_sr(pma_checker_ppn_data_barrier_7_io_x_sr),
    .io_x_pw(pma_checker_ppn_data_barrier_7_io_x_pw),
    .io_x_px(pma_checker_ppn_data_barrier_7_io_x_px),
    .io_x_pr(pma_checker_ppn_data_barrier_7_io_x_pr),
    .io_x_ppp(pma_checker_ppn_data_barrier_7_io_x_ppp),
    .io_x_pal(pma_checker_ppn_data_barrier_7_io_x_pal),
    .io_x_paa(pma_checker_ppn_data_barrier_7_io_x_paa),
    .io_x_eff(pma_checker_ppn_data_barrier_7_io_x_eff),
    .io_x_c(pma_checker_ppn_data_barrier_7_io_x_c),
    .io_y_ppn(pma_checker_ppn_data_barrier_7_io_y_ppn),
    .io_y_u(pma_checker_ppn_data_barrier_7_io_y_u),
    .io_y_ae(pma_checker_ppn_data_barrier_7_io_y_ae),
    .io_y_sw(pma_checker_ppn_data_barrier_7_io_y_sw),
    .io_y_sx(pma_checker_ppn_data_barrier_7_io_y_sx),
    .io_y_sr(pma_checker_ppn_data_barrier_7_io_y_sr),
    .io_y_pw(pma_checker_ppn_data_barrier_7_io_y_pw),
    .io_y_px(pma_checker_ppn_data_barrier_7_io_y_px),
    .io_y_pr(pma_checker_ppn_data_barrier_7_io_y_pr),
    .io_y_ppp(pma_checker_ppn_data_barrier_7_io_y_ppp),
    .io_y_pal(pma_checker_ppn_data_barrier_7_io_y_pal),
    .io_y_paa(pma_checker_ppn_data_barrier_7_io_y_paa),
    .io_y_eff(pma_checker_ppn_data_barrier_7_io_y_eff),
    .io_y_c(pma_checker_ppn_data_barrier_7_io_y_c)
  );
  OptimizationBarrier pma_checker_ppn_data_barrier_8 ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_ppn_data_barrier_8_io_x_ppn),
    .io_x_u(pma_checker_ppn_data_barrier_8_io_x_u),
    .io_x_ae(pma_checker_ppn_data_barrier_8_io_x_ae),
    .io_x_sw(pma_checker_ppn_data_barrier_8_io_x_sw),
    .io_x_sx(pma_checker_ppn_data_barrier_8_io_x_sx),
    .io_x_sr(pma_checker_ppn_data_barrier_8_io_x_sr),
    .io_x_pw(pma_checker_ppn_data_barrier_8_io_x_pw),
    .io_x_px(pma_checker_ppn_data_barrier_8_io_x_px),
    .io_x_pr(pma_checker_ppn_data_barrier_8_io_x_pr),
    .io_x_ppp(pma_checker_ppn_data_barrier_8_io_x_ppp),
    .io_x_pal(pma_checker_ppn_data_barrier_8_io_x_pal),
    .io_x_paa(pma_checker_ppn_data_barrier_8_io_x_paa),
    .io_x_eff(pma_checker_ppn_data_barrier_8_io_x_eff),
    .io_x_c(pma_checker_ppn_data_barrier_8_io_x_c),
    .io_y_ppn(pma_checker_ppn_data_barrier_8_io_y_ppn),
    .io_y_u(pma_checker_ppn_data_barrier_8_io_y_u),
    .io_y_ae(pma_checker_ppn_data_barrier_8_io_y_ae),
    .io_y_sw(pma_checker_ppn_data_barrier_8_io_y_sw),
    .io_y_sx(pma_checker_ppn_data_barrier_8_io_y_sx),
    .io_y_sr(pma_checker_ppn_data_barrier_8_io_y_sr),
    .io_y_pw(pma_checker_ppn_data_barrier_8_io_y_pw),
    .io_y_px(pma_checker_ppn_data_barrier_8_io_y_px),
    .io_y_pr(pma_checker_ppn_data_barrier_8_io_y_pr),
    .io_y_ppp(pma_checker_ppn_data_barrier_8_io_y_ppp),
    .io_y_pal(pma_checker_ppn_data_barrier_8_io_y_pal),
    .io_y_paa(pma_checker_ppn_data_barrier_8_io_y_paa),
    .io_y_eff(pma_checker_ppn_data_barrier_8_io_y_eff),
    .io_y_c(pma_checker_ppn_data_barrier_8_io_y_c)
  );
  OptimizationBarrier pma_checker_ppn_data_barrier_9 ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_ppn_data_barrier_9_io_x_ppn),
    .io_x_u(pma_checker_ppn_data_barrier_9_io_x_u),
    .io_x_ae(pma_checker_ppn_data_barrier_9_io_x_ae),
    .io_x_sw(pma_checker_ppn_data_barrier_9_io_x_sw),
    .io_x_sx(pma_checker_ppn_data_barrier_9_io_x_sx),
    .io_x_sr(pma_checker_ppn_data_barrier_9_io_x_sr),
    .io_x_pw(pma_checker_ppn_data_barrier_9_io_x_pw),
    .io_x_px(pma_checker_ppn_data_barrier_9_io_x_px),
    .io_x_pr(pma_checker_ppn_data_barrier_9_io_x_pr),
    .io_x_ppp(pma_checker_ppn_data_barrier_9_io_x_ppp),
    .io_x_pal(pma_checker_ppn_data_barrier_9_io_x_pal),
    .io_x_paa(pma_checker_ppn_data_barrier_9_io_x_paa),
    .io_x_eff(pma_checker_ppn_data_barrier_9_io_x_eff),
    .io_x_c(pma_checker_ppn_data_barrier_9_io_x_c),
    .io_y_ppn(pma_checker_ppn_data_barrier_9_io_y_ppn),
    .io_y_u(pma_checker_ppn_data_barrier_9_io_y_u),
    .io_y_ae(pma_checker_ppn_data_barrier_9_io_y_ae),
    .io_y_sw(pma_checker_ppn_data_barrier_9_io_y_sw),
    .io_y_sx(pma_checker_ppn_data_barrier_9_io_y_sx),
    .io_y_sr(pma_checker_ppn_data_barrier_9_io_y_sr),
    .io_y_pw(pma_checker_ppn_data_barrier_9_io_y_pw),
    .io_y_px(pma_checker_ppn_data_barrier_9_io_y_px),
    .io_y_pr(pma_checker_ppn_data_barrier_9_io_y_pr),
    .io_y_ppp(pma_checker_ppn_data_barrier_9_io_y_ppp),
    .io_y_pal(pma_checker_ppn_data_barrier_9_io_y_pal),
    .io_y_paa(pma_checker_ppn_data_barrier_9_io_y_paa),
    .io_y_eff(pma_checker_ppn_data_barrier_9_io_y_eff),
    .io_y_c(pma_checker_ppn_data_barrier_9_io_y_c)
  );
  OptimizationBarrier pma_checker_ppn_data_barrier_10 ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_ppn_data_barrier_10_io_x_ppn),
    .io_x_u(pma_checker_ppn_data_barrier_10_io_x_u),
    .io_x_ae(pma_checker_ppn_data_barrier_10_io_x_ae),
    .io_x_sw(pma_checker_ppn_data_barrier_10_io_x_sw),
    .io_x_sx(pma_checker_ppn_data_barrier_10_io_x_sx),
    .io_x_sr(pma_checker_ppn_data_barrier_10_io_x_sr),
    .io_x_pw(pma_checker_ppn_data_barrier_10_io_x_pw),
    .io_x_px(pma_checker_ppn_data_barrier_10_io_x_px),
    .io_x_pr(pma_checker_ppn_data_barrier_10_io_x_pr),
    .io_x_ppp(pma_checker_ppn_data_barrier_10_io_x_ppp),
    .io_x_pal(pma_checker_ppn_data_barrier_10_io_x_pal),
    .io_x_paa(pma_checker_ppn_data_barrier_10_io_x_paa),
    .io_x_eff(pma_checker_ppn_data_barrier_10_io_x_eff),
    .io_x_c(pma_checker_ppn_data_barrier_10_io_x_c),
    .io_y_ppn(pma_checker_ppn_data_barrier_10_io_y_ppn),
    .io_y_u(pma_checker_ppn_data_barrier_10_io_y_u),
    .io_y_ae(pma_checker_ppn_data_barrier_10_io_y_ae),
    .io_y_sw(pma_checker_ppn_data_barrier_10_io_y_sw),
    .io_y_sx(pma_checker_ppn_data_barrier_10_io_y_sx),
    .io_y_sr(pma_checker_ppn_data_barrier_10_io_y_sr),
    .io_y_pw(pma_checker_ppn_data_barrier_10_io_y_pw),
    .io_y_px(pma_checker_ppn_data_barrier_10_io_y_px),
    .io_y_pr(pma_checker_ppn_data_barrier_10_io_y_pr),
    .io_y_ppp(pma_checker_ppn_data_barrier_10_io_y_ppp),
    .io_y_pal(pma_checker_ppn_data_barrier_10_io_y_pal),
    .io_y_paa(pma_checker_ppn_data_barrier_10_io_y_paa),
    .io_y_eff(pma_checker_ppn_data_barrier_10_io_y_eff),
    .io_y_c(pma_checker_ppn_data_barrier_10_io_y_c)
  );
  OptimizationBarrier pma_checker_ppn_data_barrier_11 ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_ppn_data_barrier_11_io_x_ppn),
    .io_x_u(pma_checker_ppn_data_barrier_11_io_x_u),
    .io_x_ae(pma_checker_ppn_data_barrier_11_io_x_ae),
    .io_x_sw(pma_checker_ppn_data_barrier_11_io_x_sw),
    .io_x_sx(pma_checker_ppn_data_barrier_11_io_x_sx),
    .io_x_sr(pma_checker_ppn_data_barrier_11_io_x_sr),
    .io_x_pw(pma_checker_ppn_data_barrier_11_io_x_pw),
    .io_x_px(pma_checker_ppn_data_barrier_11_io_x_px),
    .io_x_pr(pma_checker_ppn_data_barrier_11_io_x_pr),
    .io_x_ppp(pma_checker_ppn_data_barrier_11_io_x_ppp),
    .io_x_pal(pma_checker_ppn_data_barrier_11_io_x_pal),
    .io_x_paa(pma_checker_ppn_data_barrier_11_io_x_paa),
    .io_x_eff(pma_checker_ppn_data_barrier_11_io_x_eff),
    .io_x_c(pma_checker_ppn_data_barrier_11_io_x_c),
    .io_y_ppn(pma_checker_ppn_data_barrier_11_io_y_ppn),
    .io_y_u(pma_checker_ppn_data_barrier_11_io_y_u),
    .io_y_ae(pma_checker_ppn_data_barrier_11_io_y_ae),
    .io_y_sw(pma_checker_ppn_data_barrier_11_io_y_sw),
    .io_y_sx(pma_checker_ppn_data_barrier_11_io_y_sx),
    .io_y_sr(pma_checker_ppn_data_barrier_11_io_y_sr),
    .io_y_pw(pma_checker_ppn_data_barrier_11_io_y_pw),
    .io_y_px(pma_checker_ppn_data_barrier_11_io_y_px),
    .io_y_pr(pma_checker_ppn_data_barrier_11_io_y_pr),
    .io_y_ppp(pma_checker_ppn_data_barrier_11_io_y_ppp),
    .io_y_pal(pma_checker_ppn_data_barrier_11_io_y_pal),
    .io_y_paa(pma_checker_ppn_data_barrier_11_io_y_paa),
    .io_y_eff(pma_checker_ppn_data_barrier_11_io_y_eff),
    .io_y_c(pma_checker_ppn_data_barrier_11_io_y_c)
  );
  OptimizationBarrier pma_checker_ppn_data_barrier_12 ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_ppn_data_barrier_12_io_x_ppn),
    .io_x_u(pma_checker_ppn_data_barrier_12_io_x_u),
    .io_x_ae(pma_checker_ppn_data_barrier_12_io_x_ae),
    .io_x_sw(pma_checker_ppn_data_barrier_12_io_x_sw),
    .io_x_sx(pma_checker_ppn_data_barrier_12_io_x_sx),
    .io_x_sr(pma_checker_ppn_data_barrier_12_io_x_sr),
    .io_x_pw(pma_checker_ppn_data_barrier_12_io_x_pw),
    .io_x_px(pma_checker_ppn_data_barrier_12_io_x_px),
    .io_x_pr(pma_checker_ppn_data_barrier_12_io_x_pr),
    .io_x_ppp(pma_checker_ppn_data_barrier_12_io_x_ppp),
    .io_x_pal(pma_checker_ppn_data_barrier_12_io_x_pal),
    .io_x_paa(pma_checker_ppn_data_barrier_12_io_x_paa),
    .io_x_eff(pma_checker_ppn_data_barrier_12_io_x_eff),
    .io_x_c(pma_checker_ppn_data_barrier_12_io_x_c),
    .io_y_ppn(pma_checker_ppn_data_barrier_12_io_y_ppn),
    .io_y_u(pma_checker_ppn_data_barrier_12_io_y_u),
    .io_y_ae(pma_checker_ppn_data_barrier_12_io_y_ae),
    .io_y_sw(pma_checker_ppn_data_barrier_12_io_y_sw),
    .io_y_sx(pma_checker_ppn_data_barrier_12_io_y_sx),
    .io_y_sr(pma_checker_ppn_data_barrier_12_io_y_sr),
    .io_y_pw(pma_checker_ppn_data_barrier_12_io_y_pw),
    .io_y_px(pma_checker_ppn_data_barrier_12_io_y_px),
    .io_y_pr(pma_checker_ppn_data_barrier_12_io_y_pr),
    .io_y_ppp(pma_checker_ppn_data_barrier_12_io_y_ppp),
    .io_y_pal(pma_checker_ppn_data_barrier_12_io_y_pal),
    .io_y_paa(pma_checker_ppn_data_barrier_12_io_y_paa),
    .io_y_eff(pma_checker_ppn_data_barrier_12_io_y_eff),
    .io_y_c(pma_checker_ppn_data_barrier_12_io_y_c)
  );
  OptimizationBarrier pma_checker_entries_barrier ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_entries_barrier_io_x_ppn),
    .io_x_u(pma_checker_entries_barrier_io_x_u),
    .io_x_ae(pma_checker_entries_barrier_io_x_ae),
    .io_x_sw(pma_checker_entries_barrier_io_x_sw),
    .io_x_sx(pma_checker_entries_barrier_io_x_sx),
    .io_x_sr(pma_checker_entries_barrier_io_x_sr),
    .io_x_pw(pma_checker_entries_barrier_io_x_pw),
    .io_x_px(pma_checker_entries_barrier_io_x_px),
    .io_x_pr(pma_checker_entries_barrier_io_x_pr),
    .io_x_ppp(pma_checker_entries_barrier_io_x_ppp),
    .io_x_pal(pma_checker_entries_barrier_io_x_pal),
    .io_x_paa(pma_checker_entries_barrier_io_x_paa),
    .io_x_eff(pma_checker_entries_barrier_io_x_eff),
    .io_x_c(pma_checker_entries_barrier_io_x_c),
    .io_y_ppn(pma_checker_entries_barrier_io_y_ppn),
    .io_y_u(pma_checker_entries_barrier_io_y_u),
    .io_y_ae(pma_checker_entries_barrier_io_y_ae),
    .io_y_sw(pma_checker_entries_barrier_io_y_sw),
    .io_y_sx(pma_checker_entries_barrier_io_y_sx),
    .io_y_sr(pma_checker_entries_barrier_io_y_sr),
    .io_y_pw(pma_checker_entries_barrier_io_y_pw),
    .io_y_px(pma_checker_entries_barrier_io_y_px),
    .io_y_pr(pma_checker_entries_barrier_io_y_pr),
    .io_y_ppp(pma_checker_entries_barrier_io_y_ppp),
    .io_y_pal(pma_checker_entries_barrier_io_y_pal),
    .io_y_paa(pma_checker_entries_barrier_io_y_paa),
    .io_y_eff(pma_checker_entries_barrier_io_y_eff),
    .io_y_c(pma_checker_entries_barrier_io_y_c)
  );
  OptimizationBarrier pma_checker_entries_barrier_1 ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_entries_barrier_1_io_x_ppn),
    .io_x_u(pma_checker_entries_barrier_1_io_x_u),
    .io_x_ae(pma_checker_entries_barrier_1_io_x_ae),
    .io_x_sw(pma_checker_entries_barrier_1_io_x_sw),
    .io_x_sx(pma_checker_entries_barrier_1_io_x_sx),
    .io_x_sr(pma_checker_entries_barrier_1_io_x_sr),
    .io_x_pw(pma_checker_entries_barrier_1_io_x_pw),
    .io_x_px(pma_checker_entries_barrier_1_io_x_px),
    .io_x_pr(pma_checker_entries_barrier_1_io_x_pr),
    .io_x_ppp(pma_checker_entries_barrier_1_io_x_ppp),
    .io_x_pal(pma_checker_entries_barrier_1_io_x_pal),
    .io_x_paa(pma_checker_entries_barrier_1_io_x_paa),
    .io_x_eff(pma_checker_entries_barrier_1_io_x_eff),
    .io_x_c(pma_checker_entries_barrier_1_io_x_c),
    .io_y_ppn(pma_checker_entries_barrier_1_io_y_ppn),
    .io_y_u(pma_checker_entries_barrier_1_io_y_u),
    .io_y_ae(pma_checker_entries_barrier_1_io_y_ae),
    .io_y_sw(pma_checker_entries_barrier_1_io_y_sw),
    .io_y_sx(pma_checker_entries_barrier_1_io_y_sx),
    .io_y_sr(pma_checker_entries_barrier_1_io_y_sr),
    .io_y_pw(pma_checker_entries_barrier_1_io_y_pw),
    .io_y_px(pma_checker_entries_barrier_1_io_y_px),
    .io_y_pr(pma_checker_entries_barrier_1_io_y_pr),
    .io_y_ppp(pma_checker_entries_barrier_1_io_y_ppp),
    .io_y_pal(pma_checker_entries_barrier_1_io_y_pal),
    .io_y_paa(pma_checker_entries_barrier_1_io_y_paa),
    .io_y_eff(pma_checker_entries_barrier_1_io_y_eff),
    .io_y_c(pma_checker_entries_barrier_1_io_y_c)
  );
  OptimizationBarrier pma_checker_entries_barrier_2 ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_entries_barrier_2_io_x_ppn),
    .io_x_u(pma_checker_entries_barrier_2_io_x_u),
    .io_x_ae(pma_checker_entries_barrier_2_io_x_ae),
    .io_x_sw(pma_checker_entries_barrier_2_io_x_sw),
    .io_x_sx(pma_checker_entries_barrier_2_io_x_sx),
    .io_x_sr(pma_checker_entries_barrier_2_io_x_sr),
    .io_x_pw(pma_checker_entries_barrier_2_io_x_pw),
    .io_x_px(pma_checker_entries_barrier_2_io_x_px),
    .io_x_pr(pma_checker_entries_barrier_2_io_x_pr),
    .io_x_ppp(pma_checker_entries_barrier_2_io_x_ppp),
    .io_x_pal(pma_checker_entries_barrier_2_io_x_pal),
    .io_x_paa(pma_checker_entries_barrier_2_io_x_paa),
    .io_x_eff(pma_checker_entries_barrier_2_io_x_eff),
    .io_x_c(pma_checker_entries_barrier_2_io_x_c),
    .io_y_ppn(pma_checker_entries_barrier_2_io_y_ppn),
    .io_y_u(pma_checker_entries_barrier_2_io_y_u),
    .io_y_ae(pma_checker_entries_barrier_2_io_y_ae),
    .io_y_sw(pma_checker_entries_barrier_2_io_y_sw),
    .io_y_sx(pma_checker_entries_barrier_2_io_y_sx),
    .io_y_sr(pma_checker_entries_barrier_2_io_y_sr),
    .io_y_pw(pma_checker_entries_barrier_2_io_y_pw),
    .io_y_px(pma_checker_entries_barrier_2_io_y_px),
    .io_y_pr(pma_checker_entries_barrier_2_io_y_pr),
    .io_y_ppp(pma_checker_entries_barrier_2_io_y_ppp),
    .io_y_pal(pma_checker_entries_barrier_2_io_y_pal),
    .io_y_paa(pma_checker_entries_barrier_2_io_y_paa),
    .io_y_eff(pma_checker_entries_barrier_2_io_y_eff),
    .io_y_c(pma_checker_entries_barrier_2_io_y_c)
  );
  OptimizationBarrier pma_checker_entries_barrier_3 ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_entries_barrier_3_io_x_ppn),
    .io_x_u(pma_checker_entries_barrier_3_io_x_u),
    .io_x_ae(pma_checker_entries_barrier_3_io_x_ae),
    .io_x_sw(pma_checker_entries_barrier_3_io_x_sw),
    .io_x_sx(pma_checker_entries_barrier_3_io_x_sx),
    .io_x_sr(pma_checker_entries_barrier_3_io_x_sr),
    .io_x_pw(pma_checker_entries_barrier_3_io_x_pw),
    .io_x_px(pma_checker_entries_barrier_3_io_x_px),
    .io_x_pr(pma_checker_entries_barrier_3_io_x_pr),
    .io_x_ppp(pma_checker_entries_barrier_3_io_x_ppp),
    .io_x_pal(pma_checker_entries_barrier_3_io_x_pal),
    .io_x_paa(pma_checker_entries_barrier_3_io_x_paa),
    .io_x_eff(pma_checker_entries_barrier_3_io_x_eff),
    .io_x_c(pma_checker_entries_barrier_3_io_x_c),
    .io_y_ppn(pma_checker_entries_barrier_3_io_y_ppn),
    .io_y_u(pma_checker_entries_barrier_3_io_y_u),
    .io_y_ae(pma_checker_entries_barrier_3_io_y_ae),
    .io_y_sw(pma_checker_entries_barrier_3_io_y_sw),
    .io_y_sx(pma_checker_entries_barrier_3_io_y_sx),
    .io_y_sr(pma_checker_entries_barrier_3_io_y_sr),
    .io_y_pw(pma_checker_entries_barrier_3_io_y_pw),
    .io_y_px(pma_checker_entries_barrier_3_io_y_px),
    .io_y_pr(pma_checker_entries_barrier_3_io_y_pr),
    .io_y_ppp(pma_checker_entries_barrier_3_io_y_ppp),
    .io_y_pal(pma_checker_entries_barrier_3_io_y_pal),
    .io_y_paa(pma_checker_entries_barrier_3_io_y_paa),
    .io_y_eff(pma_checker_entries_barrier_3_io_y_eff),
    .io_y_c(pma_checker_entries_barrier_3_io_y_c)
  );
  OptimizationBarrier pma_checker_entries_barrier_4 ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_entries_barrier_4_io_x_ppn),
    .io_x_u(pma_checker_entries_barrier_4_io_x_u),
    .io_x_ae(pma_checker_entries_barrier_4_io_x_ae),
    .io_x_sw(pma_checker_entries_barrier_4_io_x_sw),
    .io_x_sx(pma_checker_entries_barrier_4_io_x_sx),
    .io_x_sr(pma_checker_entries_barrier_4_io_x_sr),
    .io_x_pw(pma_checker_entries_barrier_4_io_x_pw),
    .io_x_px(pma_checker_entries_barrier_4_io_x_px),
    .io_x_pr(pma_checker_entries_barrier_4_io_x_pr),
    .io_x_ppp(pma_checker_entries_barrier_4_io_x_ppp),
    .io_x_pal(pma_checker_entries_barrier_4_io_x_pal),
    .io_x_paa(pma_checker_entries_barrier_4_io_x_paa),
    .io_x_eff(pma_checker_entries_barrier_4_io_x_eff),
    .io_x_c(pma_checker_entries_barrier_4_io_x_c),
    .io_y_ppn(pma_checker_entries_barrier_4_io_y_ppn),
    .io_y_u(pma_checker_entries_barrier_4_io_y_u),
    .io_y_ae(pma_checker_entries_barrier_4_io_y_ae),
    .io_y_sw(pma_checker_entries_barrier_4_io_y_sw),
    .io_y_sx(pma_checker_entries_barrier_4_io_y_sx),
    .io_y_sr(pma_checker_entries_barrier_4_io_y_sr),
    .io_y_pw(pma_checker_entries_barrier_4_io_y_pw),
    .io_y_px(pma_checker_entries_barrier_4_io_y_px),
    .io_y_pr(pma_checker_entries_barrier_4_io_y_pr),
    .io_y_ppp(pma_checker_entries_barrier_4_io_y_ppp),
    .io_y_pal(pma_checker_entries_barrier_4_io_y_pal),
    .io_y_paa(pma_checker_entries_barrier_4_io_y_paa),
    .io_y_eff(pma_checker_entries_barrier_4_io_y_eff),
    .io_y_c(pma_checker_entries_barrier_4_io_y_c)
  );
  OptimizationBarrier pma_checker_entries_barrier_5 ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_entries_barrier_5_io_x_ppn),
    .io_x_u(pma_checker_entries_barrier_5_io_x_u),
    .io_x_ae(pma_checker_entries_barrier_5_io_x_ae),
    .io_x_sw(pma_checker_entries_barrier_5_io_x_sw),
    .io_x_sx(pma_checker_entries_barrier_5_io_x_sx),
    .io_x_sr(pma_checker_entries_barrier_5_io_x_sr),
    .io_x_pw(pma_checker_entries_barrier_5_io_x_pw),
    .io_x_px(pma_checker_entries_barrier_5_io_x_px),
    .io_x_pr(pma_checker_entries_barrier_5_io_x_pr),
    .io_x_ppp(pma_checker_entries_barrier_5_io_x_ppp),
    .io_x_pal(pma_checker_entries_barrier_5_io_x_pal),
    .io_x_paa(pma_checker_entries_barrier_5_io_x_paa),
    .io_x_eff(pma_checker_entries_barrier_5_io_x_eff),
    .io_x_c(pma_checker_entries_barrier_5_io_x_c),
    .io_y_ppn(pma_checker_entries_barrier_5_io_y_ppn),
    .io_y_u(pma_checker_entries_barrier_5_io_y_u),
    .io_y_ae(pma_checker_entries_barrier_5_io_y_ae),
    .io_y_sw(pma_checker_entries_barrier_5_io_y_sw),
    .io_y_sx(pma_checker_entries_barrier_5_io_y_sx),
    .io_y_sr(pma_checker_entries_barrier_5_io_y_sr),
    .io_y_pw(pma_checker_entries_barrier_5_io_y_pw),
    .io_y_px(pma_checker_entries_barrier_5_io_y_px),
    .io_y_pr(pma_checker_entries_barrier_5_io_y_pr),
    .io_y_ppp(pma_checker_entries_barrier_5_io_y_ppp),
    .io_y_pal(pma_checker_entries_barrier_5_io_y_pal),
    .io_y_paa(pma_checker_entries_barrier_5_io_y_paa),
    .io_y_eff(pma_checker_entries_barrier_5_io_y_eff),
    .io_y_c(pma_checker_entries_barrier_5_io_y_c)
  );
  OptimizationBarrier pma_checker_entries_barrier_6 ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_entries_barrier_6_io_x_ppn),
    .io_x_u(pma_checker_entries_barrier_6_io_x_u),
    .io_x_ae(pma_checker_entries_barrier_6_io_x_ae),
    .io_x_sw(pma_checker_entries_barrier_6_io_x_sw),
    .io_x_sx(pma_checker_entries_barrier_6_io_x_sx),
    .io_x_sr(pma_checker_entries_barrier_6_io_x_sr),
    .io_x_pw(pma_checker_entries_barrier_6_io_x_pw),
    .io_x_px(pma_checker_entries_barrier_6_io_x_px),
    .io_x_pr(pma_checker_entries_barrier_6_io_x_pr),
    .io_x_ppp(pma_checker_entries_barrier_6_io_x_ppp),
    .io_x_pal(pma_checker_entries_barrier_6_io_x_pal),
    .io_x_paa(pma_checker_entries_barrier_6_io_x_paa),
    .io_x_eff(pma_checker_entries_barrier_6_io_x_eff),
    .io_x_c(pma_checker_entries_barrier_6_io_x_c),
    .io_y_ppn(pma_checker_entries_barrier_6_io_y_ppn),
    .io_y_u(pma_checker_entries_barrier_6_io_y_u),
    .io_y_ae(pma_checker_entries_barrier_6_io_y_ae),
    .io_y_sw(pma_checker_entries_barrier_6_io_y_sw),
    .io_y_sx(pma_checker_entries_barrier_6_io_y_sx),
    .io_y_sr(pma_checker_entries_barrier_6_io_y_sr),
    .io_y_pw(pma_checker_entries_barrier_6_io_y_pw),
    .io_y_px(pma_checker_entries_barrier_6_io_y_px),
    .io_y_pr(pma_checker_entries_barrier_6_io_y_pr),
    .io_y_ppp(pma_checker_entries_barrier_6_io_y_ppp),
    .io_y_pal(pma_checker_entries_barrier_6_io_y_pal),
    .io_y_paa(pma_checker_entries_barrier_6_io_y_paa),
    .io_y_eff(pma_checker_entries_barrier_6_io_y_eff),
    .io_y_c(pma_checker_entries_barrier_6_io_y_c)
  );
  OptimizationBarrier pma_checker_entries_barrier_7 ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_entries_barrier_7_io_x_ppn),
    .io_x_u(pma_checker_entries_barrier_7_io_x_u),
    .io_x_ae(pma_checker_entries_barrier_7_io_x_ae),
    .io_x_sw(pma_checker_entries_barrier_7_io_x_sw),
    .io_x_sx(pma_checker_entries_barrier_7_io_x_sx),
    .io_x_sr(pma_checker_entries_barrier_7_io_x_sr),
    .io_x_pw(pma_checker_entries_barrier_7_io_x_pw),
    .io_x_px(pma_checker_entries_barrier_7_io_x_px),
    .io_x_pr(pma_checker_entries_barrier_7_io_x_pr),
    .io_x_ppp(pma_checker_entries_barrier_7_io_x_ppp),
    .io_x_pal(pma_checker_entries_barrier_7_io_x_pal),
    .io_x_paa(pma_checker_entries_barrier_7_io_x_paa),
    .io_x_eff(pma_checker_entries_barrier_7_io_x_eff),
    .io_x_c(pma_checker_entries_barrier_7_io_x_c),
    .io_y_ppn(pma_checker_entries_barrier_7_io_y_ppn),
    .io_y_u(pma_checker_entries_barrier_7_io_y_u),
    .io_y_ae(pma_checker_entries_barrier_7_io_y_ae),
    .io_y_sw(pma_checker_entries_barrier_7_io_y_sw),
    .io_y_sx(pma_checker_entries_barrier_7_io_y_sx),
    .io_y_sr(pma_checker_entries_barrier_7_io_y_sr),
    .io_y_pw(pma_checker_entries_barrier_7_io_y_pw),
    .io_y_px(pma_checker_entries_barrier_7_io_y_px),
    .io_y_pr(pma_checker_entries_barrier_7_io_y_pr),
    .io_y_ppp(pma_checker_entries_barrier_7_io_y_ppp),
    .io_y_pal(pma_checker_entries_barrier_7_io_y_pal),
    .io_y_paa(pma_checker_entries_barrier_7_io_y_paa),
    .io_y_eff(pma_checker_entries_barrier_7_io_y_eff),
    .io_y_c(pma_checker_entries_barrier_7_io_y_c)
  );
  OptimizationBarrier pma_checker_entries_barrier_8 ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_entries_barrier_8_io_x_ppn),
    .io_x_u(pma_checker_entries_barrier_8_io_x_u),
    .io_x_ae(pma_checker_entries_barrier_8_io_x_ae),
    .io_x_sw(pma_checker_entries_barrier_8_io_x_sw),
    .io_x_sx(pma_checker_entries_barrier_8_io_x_sx),
    .io_x_sr(pma_checker_entries_barrier_8_io_x_sr),
    .io_x_pw(pma_checker_entries_barrier_8_io_x_pw),
    .io_x_px(pma_checker_entries_barrier_8_io_x_px),
    .io_x_pr(pma_checker_entries_barrier_8_io_x_pr),
    .io_x_ppp(pma_checker_entries_barrier_8_io_x_ppp),
    .io_x_pal(pma_checker_entries_barrier_8_io_x_pal),
    .io_x_paa(pma_checker_entries_barrier_8_io_x_paa),
    .io_x_eff(pma_checker_entries_barrier_8_io_x_eff),
    .io_x_c(pma_checker_entries_barrier_8_io_x_c),
    .io_y_ppn(pma_checker_entries_barrier_8_io_y_ppn),
    .io_y_u(pma_checker_entries_barrier_8_io_y_u),
    .io_y_ae(pma_checker_entries_barrier_8_io_y_ae),
    .io_y_sw(pma_checker_entries_barrier_8_io_y_sw),
    .io_y_sx(pma_checker_entries_barrier_8_io_y_sx),
    .io_y_sr(pma_checker_entries_barrier_8_io_y_sr),
    .io_y_pw(pma_checker_entries_barrier_8_io_y_pw),
    .io_y_px(pma_checker_entries_barrier_8_io_y_px),
    .io_y_pr(pma_checker_entries_barrier_8_io_y_pr),
    .io_y_ppp(pma_checker_entries_barrier_8_io_y_ppp),
    .io_y_pal(pma_checker_entries_barrier_8_io_y_pal),
    .io_y_paa(pma_checker_entries_barrier_8_io_y_paa),
    .io_y_eff(pma_checker_entries_barrier_8_io_y_eff),
    .io_y_c(pma_checker_entries_barrier_8_io_y_c)
  );
  OptimizationBarrier pma_checker_entries_barrier_9 ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_entries_barrier_9_io_x_ppn),
    .io_x_u(pma_checker_entries_barrier_9_io_x_u),
    .io_x_ae(pma_checker_entries_barrier_9_io_x_ae),
    .io_x_sw(pma_checker_entries_barrier_9_io_x_sw),
    .io_x_sx(pma_checker_entries_barrier_9_io_x_sx),
    .io_x_sr(pma_checker_entries_barrier_9_io_x_sr),
    .io_x_pw(pma_checker_entries_barrier_9_io_x_pw),
    .io_x_px(pma_checker_entries_barrier_9_io_x_px),
    .io_x_pr(pma_checker_entries_barrier_9_io_x_pr),
    .io_x_ppp(pma_checker_entries_barrier_9_io_x_ppp),
    .io_x_pal(pma_checker_entries_barrier_9_io_x_pal),
    .io_x_paa(pma_checker_entries_barrier_9_io_x_paa),
    .io_x_eff(pma_checker_entries_barrier_9_io_x_eff),
    .io_x_c(pma_checker_entries_barrier_9_io_x_c),
    .io_y_ppn(pma_checker_entries_barrier_9_io_y_ppn),
    .io_y_u(pma_checker_entries_barrier_9_io_y_u),
    .io_y_ae(pma_checker_entries_barrier_9_io_y_ae),
    .io_y_sw(pma_checker_entries_barrier_9_io_y_sw),
    .io_y_sx(pma_checker_entries_barrier_9_io_y_sx),
    .io_y_sr(pma_checker_entries_barrier_9_io_y_sr),
    .io_y_pw(pma_checker_entries_barrier_9_io_y_pw),
    .io_y_px(pma_checker_entries_barrier_9_io_y_px),
    .io_y_pr(pma_checker_entries_barrier_9_io_y_pr),
    .io_y_ppp(pma_checker_entries_barrier_9_io_y_ppp),
    .io_y_pal(pma_checker_entries_barrier_9_io_y_pal),
    .io_y_paa(pma_checker_entries_barrier_9_io_y_paa),
    .io_y_eff(pma_checker_entries_barrier_9_io_y_eff),
    .io_y_c(pma_checker_entries_barrier_9_io_y_c)
  );
  OptimizationBarrier pma_checker_entries_barrier_10 ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_entries_barrier_10_io_x_ppn),
    .io_x_u(pma_checker_entries_barrier_10_io_x_u),
    .io_x_ae(pma_checker_entries_barrier_10_io_x_ae),
    .io_x_sw(pma_checker_entries_barrier_10_io_x_sw),
    .io_x_sx(pma_checker_entries_barrier_10_io_x_sx),
    .io_x_sr(pma_checker_entries_barrier_10_io_x_sr),
    .io_x_pw(pma_checker_entries_barrier_10_io_x_pw),
    .io_x_px(pma_checker_entries_barrier_10_io_x_px),
    .io_x_pr(pma_checker_entries_barrier_10_io_x_pr),
    .io_x_ppp(pma_checker_entries_barrier_10_io_x_ppp),
    .io_x_pal(pma_checker_entries_barrier_10_io_x_pal),
    .io_x_paa(pma_checker_entries_barrier_10_io_x_paa),
    .io_x_eff(pma_checker_entries_barrier_10_io_x_eff),
    .io_x_c(pma_checker_entries_barrier_10_io_x_c),
    .io_y_ppn(pma_checker_entries_barrier_10_io_y_ppn),
    .io_y_u(pma_checker_entries_barrier_10_io_y_u),
    .io_y_ae(pma_checker_entries_barrier_10_io_y_ae),
    .io_y_sw(pma_checker_entries_barrier_10_io_y_sw),
    .io_y_sx(pma_checker_entries_barrier_10_io_y_sx),
    .io_y_sr(pma_checker_entries_barrier_10_io_y_sr),
    .io_y_pw(pma_checker_entries_barrier_10_io_y_pw),
    .io_y_px(pma_checker_entries_barrier_10_io_y_px),
    .io_y_pr(pma_checker_entries_barrier_10_io_y_pr),
    .io_y_ppp(pma_checker_entries_barrier_10_io_y_ppp),
    .io_y_pal(pma_checker_entries_barrier_10_io_y_pal),
    .io_y_paa(pma_checker_entries_barrier_10_io_y_paa),
    .io_y_eff(pma_checker_entries_barrier_10_io_y_eff),
    .io_y_c(pma_checker_entries_barrier_10_io_y_c)
  );
  OptimizationBarrier pma_checker_entries_barrier_11 ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_entries_barrier_11_io_x_ppn),
    .io_x_u(pma_checker_entries_barrier_11_io_x_u),
    .io_x_ae(pma_checker_entries_barrier_11_io_x_ae),
    .io_x_sw(pma_checker_entries_barrier_11_io_x_sw),
    .io_x_sx(pma_checker_entries_barrier_11_io_x_sx),
    .io_x_sr(pma_checker_entries_barrier_11_io_x_sr),
    .io_x_pw(pma_checker_entries_barrier_11_io_x_pw),
    .io_x_px(pma_checker_entries_barrier_11_io_x_px),
    .io_x_pr(pma_checker_entries_barrier_11_io_x_pr),
    .io_x_ppp(pma_checker_entries_barrier_11_io_x_ppp),
    .io_x_pal(pma_checker_entries_barrier_11_io_x_pal),
    .io_x_paa(pma_checker_entries_barrier_11_io_x_paa),
    .io_x_eff(pma_checker_entries_barrier_11_io_x_eff),
    .io_x_c(pma_checker_entries_barrier_11_io_x_c),
    .io_y_ppn(pma_checker_entries_barrier_11_io_y_ppn),
    .io_y_u(pma_checker_entries_barrier_11_io_y_u),
    .io_y_ae(pma_checker_entries_barrier_11_io_y_ae),
    .io_y_sw(pma_checker_entries_barrier_11_io_y_sw),
    .io_y_sx(pma_checker_entries_barrier_11_io_y_sx),
    .io_y_sr(pma_checker_entries_barrier_11_io_y_sr),
    .io_y_pw(pma_checker_entries_barrier_11_io_y_pw),
    .io_y_px(pma_checker_entries_barrier_11_io_y_px),
    .io_y_pr(pma_checker_entries_barrier_11_io_y_pr),
    .io_y_ppp(pma_checker_entries_barrier_11_io_y_ppp),
    .io_y_pal(pma_checker_entries_barrier_11_io_y_pal),
    .io_y_paa(pma_checker_entries_barrier_11_io_y_paa),
    .io_y_eff(pma_checker_entries_barrier_11_io_y_eff),
    .io_y_c(pma_checker_entries_barrier_11_io_y_c)
  );
  OptimizationBarrier pma_checker_entries_barrier_12 ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_entries_barrier_12_io_x_ppn),
    .io_x_u(pma_checker_entries_barrier_12_io_x_u),
    .io_x_ae(pma_checker_entries_barrier_12_io_x_ae),
    .io_x_sw(pma_checker_entries_barrier_12_io_x_sw),
    .io_x_sx(pma_checker_entries_barrier_12_io_x_sx),
    .io_x_sr(pma_checker_entries_barrier_12_io_x_sr),
    .io_x_pw(pma_checker_entries_barrier_12_io_x_pw),
    .io_x_px(pma_checker_entries_barrier_12_io_x_px),
    .io_x_pr(pma_checker_entries_barrier_12_io_x_pr),
    .io_x_ppp(pma_checker_entries_barrier_12_io_x_ppp),
    .io_x_pal(pma_checker_entries_barrier_12_io_x_pal),
    .io_x_paa(pma_checker_entries_barrier_12_io_x_paa),
    .io_x_eff(pma_checker_entries_barrier_12_io_x_eff),
    .io_x_c(pma_checker_entries_barrier_12_io_x_c),
    .io_y_ppn(pma_checker_entries_barrier_12_io_y_ppn),
    .io_y_u(pma_checker_entries_barrier_12_io_y_u),
    .io_y_ae(pma_checker_entries_barrier_12_io_y_ae),
    .io_y_sw(pma_checker_entries_barrier_12_io_y_sw),
    .io_y_sx(pma_checker_entries_barrier_12_io_y_sx),
    .io_y_sr(pma_checker_entries_barrier_12_io_y_sr),
    .io_y_pw(pma_checker_entries_barrier_12_io_y_pw),
    .io_y_px(pma_checker_entries_barrier_12_io_y_px),
    .io_y_pr(pma_checker_entries_barrier_12_io_y_pr),
    .io_y_ppp(pma_checker_entries_barrier_12_io_y_ppp),
    .io_y_pal(pma_checker_entries_barrier_12_io_y_pal),
    .io_y_paa(pma_checker_entries_barrier_12_io_y_paa),
    .io_y_eff(pma_checker_entries_barrier_12_io_y_eff),
    .io_y_c(pma_checker_entries_barrier_12_io_y_c)
  );
  OptimizationBarrier pma_checker_normal_entries_barrier ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_normal_entries_barrier_io_x_ppn),
    .io_x_u(pma_checker_normal_entries_barrier_io_x_u),
    .io_x_ae(pma_checker_normal_entries_barrier_io_x_ae),
    .io_x_sw(pma_checker_normal_entries_barrier_io_x_sw),
    .io_x_sx(pma_checker_normal_entries_barrier_io_x_sx),
    .io_x_sr(pma_checker_normal_entries_barrier_io_x_sr),
    .io_x_pw(pma_checker_normal_entries_barrier_io_x_pw),
    .io_x_px(pma_checker_normal_entries_barrier_io_x_px),
    .io_x_pr(pma_checker_normal_entries_barrier_io_x_pr),
    .io_x_ppp(pma_checker_normal_entries_barrier_io_x_ppp),
    .io_x_pal(pma_checker_normal_entries_barrier_io_x_pal),
    .io_x_paa(pma_checker_normal_entries_barrier_io_x_paa),
    .io_x_eff(pma_checker_normal_entries_barrier_io_x_eff),
    .io_x_c(pma_checker_normal_entries_barrier_io_x_c),
    .io_y_ppn(pma_checker_normal_entries_barrier_io_y_ppn),
    .io_y_u(pma_checker_normal_entries_barrier_io_y_u),
    .io_y_ae(pma_checker_normal_entries_barrier_io_y_ae),
    .io_y_sw(pma_checker_normal_entries_barrier_io_y_sw),
    .io_y_sx(pma_checker_normal_entries_barrier_io_y_sx),
    .io_y_sr(pma_checker_normal_entries_barrier_io_y_sr),
    .io_y_pw(pma_checker_normal_entries_barrier_io_y_pw),
    .io_y_px(pma_checker_normal_entries_barrier_io_y_px),
    .io_y_pr(pma_checker_normal_entries_barrier_io_y_pr),
    .io_y_ppp(pma_checker_normal_entries_barrier_io_y_ppp),
    .io_y_pal(pma_checker_normal_entries_barrier_io_y_pal),
    .io_y_paa(pma_checker_normal_entries_barrier_io_y_paa),
    .io_y_eff(pma_checker_normal_entries_barrier_io_y_eff),
    .io_y_c(pma_checker_normal_entries_barrier_io_y_c)
  );
  OptimizationBarrier pma_checker_normal_entries_barrier_1 ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_normal_entries_barrier_1_io_x_ppn),
    .io_x_u(pma_checker_normal_entries_barrier_1_io_x_u),
    .io_x_ae(pma_checker_normal_entries_barrier_1_io_x_ae),
    .io_x_sw(pma_checker_normal_entries_barrier_1_io_x_sw),
    .io_x_sx(pma_checker_normal_entries_barrier_1_io_x_sx),
    .io_x_sr(pma_checker_normal_entries_barrier_1_io_x_sr),
    .io_x_pw(pma_checker_normal_entries_barrier_1_io_x_pw),
    .io_x_px(pma_checker_normal_entries_barrier_1_io_x_px),
    .io_x_pr(pma_checker_normal_entries_barrier_1_io_x_pr),
    .io_x_ppp(pma_checker_normal_entries_barrier_1_io_x_ppp),
    .io_x_pal(pma_checker_normal_entries_barrier_1_io_x_pal),
    .io_x_paa(pma_checker_normal_entries_barrier_1_io_x_paa),
    .io_x_eff(pma_checker_normal_entries_barrier_1_io_x_eff),
    .io_x_c(pma_checker_normal_entries_barrier_1_io_x_c),
    .io_y_ppn(pma_checker_normal_entries_barrier_1_io_y_ppn),
    .io_y_u(pma_checker_normal_entries_barrier_1_io_y_u),
    .io_y_ae(pma_checker_normal_entries_barrier_1_io_y_ae),
    .io_y_sw(pma_checker_normal_entries_barrier_1_io_y_sw),
    .io_y_sx(pma_checker_normal_entries_barrier_1_io_y_sx),
    .io_y_sr(pma_checker_normal_entries_barrier_1_io_y_sr),
    .io_y_pw(pma_checker_normal_entries_barrier_1_io_y_pw),
    .io_y_px(pma_checker_normal_entries_barrier_1_io_y_px),
    .io_y_pr(pma_checker_normal_entries_barrier_1_io_y_pr),
    .io_y_ppp(pma_checker_normal_entries_barrier_1_io_y_ppp),
    .io_y_pal(pma_checker_normal_entries_barrier_1_io_y_pal),
    .io_y_paa(pma_checker_normal_entries_barrier_1_io_y_paa),
    .io_y_eff(pma_checker_normal_entries_barrier_1_io_y_eff),
    .io_y_c(pma_checker_normal_entries_barrier_1_io_y_c)
  );
  OptimizationBarrier pma_checker_normal_entries_barrier_2 ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_normal_entries_barrier_2_io_x_ppn),
    .io_x_u(pma_checker_normal_entries_barrier_2_io_x_u),
    .io_x_ae(pma_checker_normal_entries_barrier_2_io_x_ae),
    .io_x_sw(pma_checker_normal_entries_barrier_2_io_x_sw),
    .io_x_sx(pma_checker_normal_entries_barrier_2_io_x_sx),
    .io_x_sr(pma_checker_normal_entries_barrier_2_io_x_sr),
    .io_x_pw(pma_checker_normal_entries_barrier_2_io_x_pw),
    .io_x_px(pma_checker_normal_entries_barrier_2_io_x_px),
    .io_x_pr(pma_checker_normal_entries_barrier_2_io_x_pr),
    .io_x_ppp(pma_checker_normal_entries_barrier_2_io_x_ppp),
    .io_x_pal(pma_checker_normal_entries_barrier_2_io_x_pal),
    .io_x_paa(pma_checker_normal_entries_barrier_2_io_x_paa),
    .io_x_eff(pma_checker_normal_entries_barrier_2_io_x_eff),
    .io_x_c(pma_checker_normal_entries_barrier_2_io_x_c),
    .io_y_ppn(pma_checker_normal_entries_barrier_2_io_y_ppn),
    .io_y_u(pma_checker_normal_entries_barrier_2_io_y_u),
    .io_y_ae(pma_checker_normal_entries_barrier_2_io_y_ae),
    .io_y_sw(pma_checker_normal_entries_barrier_2_io_y_sw),
    .io_y_sx(pma_checker_normal_entries_barrier_2_io_y_sx),
    .io_y_sr(pma_checker_normal_entries_barrier_2_io_y_sr),
    .io_y_pw(pma_checker_normal_entries_barrier_2_io_y_pw),
    .io_y_px(pma_checker_normal_entries_barrier_2_io_y_px),
    .io_y_pr(pma_checker_normal_entries_barrier_2_io_y_pr),
    .io_y_ppp(pma_checker_normal_entries_barrier_2_io_y_ppp),
    .io_y_pal(pma_checker_normal_entries_barrier_2_io_y_pal),
    .io_y_paa(pma_checker_normal_entries_barrier_2_io_y_paa),
    .io_y_eff(pma_checker_normal_entries_barrier_2_io_y_eff),
    .io_y_c(pma_checker_normal_entries_barrier_2_io_y_c)
  );
  OptimizationBarrier pma_checker_normal_entries_barrier_3 ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_normal_entries_barrier_3_io_x_ppn),
    .io_x_u(pma_checker_normal_entries_barrier_3_io_x_u),
    .io_x_ae(pma_checker_normal_entries_barrier_3_io_x_ae),
    .io_x_sw(pma_checker_normal_entries_barrier_3_io_x_sw),
    .io_x_sx(pma_checker_normal_entries_barrier_3_io_x_sx),
    .io_x_sr(pma_checker_normal_entries_barrier_3_io_x_sr),
    .io_x_pw(pma_checker_normal_entries_barrier_3_io_x_pw),
    .io_x_px(pma_checker_normal_entries_barrier_3_io_x_px),
    .io_x_pr(pma_checker_normal_entries_barrier_3_io_x_pr),
    .io_x_ppp(pma_checker_normal_entries_barrier_3_io_x_ppp),
    .io_x_pal(pma_checker_normal_entries_barrier_3_io_x_pal),
    .io_x_paa(pma_checker_normal_entries_barrier_3_io_x_paa),
    .io_x_eff(pma_checker_normal_entries_barrier_3_io_x_eff),
    .io_x_c(pma_checker_normal_entries_barrier_3_io_x_c),
    .io_y_ppn(pma_checker_normal_entries_barrier_3_io_y_ppn),
    .io_y_u(pma_checker_normal_entries_barrier_3_io_y_u),
    .io_y_ae(pma_checker_normal_entries_barrier_3_io_y_ae),
    .io_y_sw(pma_checker_normal_entries_barrier_3_io_y_sw),
    .io_y_sx(pma_checker_normal_entries_barrier_3_io_y_sx),
    .io_y_sr(pma_checker_normal_entries_barrier_3_io_y_sr),
    .io_y_pw(pma_checker_normal_entries_barrier_3_io_y_pw),
    .io_y_px(pma_checker_normal_entries_barrier_3_io_y_px),
    .io_y_pr(pma_checker_normal_entries_barrier_3_io_y_pr),
    .io_y_ppp(pma_checker_normal_entries_barrier_3_io_y_ppp),
    .io_y_pal(pma_checker_normal_entries_barrier_3_io_y_pal),
    .io_y_paa(pma_checker_normal_entries_barrier_3_io_y_paa),
    .io_y_eff(pma_checker_normal_entries_barrier_3_io_y_eff),
    .io_y_c(pma_checker_normal_entries_barrier_3_io_y_c)
  );
  OptimizationBarrier pma_checker_normal_entries_barrier_4 ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_normal_entries_barrier_4_io_x_ppn),
    .io_x_u(pma_checker_normal_entries_barrier_4_io_x_u),
    .io_x_ae(pma_checker_normal_entries_barrier_4_io_x_ae),
    .io_x_sw(pma_checker_normal_entries_barrier_4_io_x_sw),
    .io_x_sx(pma_checker_normal_entries_barrier_4_io_x_sx),
    .io_x_sr(pma_checker_normal_entries_barrier_4_io_x_sr),
    .io_x_pw(pma_checker_normal_entries_barrier_4_io_x_pw),
    .io_x_px(pma_checker_normal_entries_barrier_4_io_x_px),
    .io_x_pr(pma_checker_normal_entries_barrier_4_io_x_pr),
    .io_x_ppp(pma_checker_normal_entries_barrier_4_io_x_ppp),
    .io_x_pal(pma_checker_normal_entries_barrier_4_io_x_pal),
    .io_x_paa(pma_checker_normal_entries_barrier_4_io_x_paa),
    .io_x_eff(pma_checker_normal_entries_barrier_4_io_x_eff),
    .io_x_c(pma_checker_normal_entries_barrier_4_io_x_c),
    .io_y_ppn(pma_checker_normal_entries_barrier_4_io_y_ppn),
    .io_y_u(pma_checker_normal_entries_barrier_4_io_y_u),
    .io_y_ae(pma_checker_normal_entries_barrier_4_io_y_ae),
    .io_y_sw(pma_checker_normal_entries_barrier_4_io_y_sw),
    .io_y_sx(pma_checker_normal_entries_barrier_4_io_y_sx),
    .io_y_sr(pma_checker_normal_entries_barrier_4_io_y_sr),
    .io_y_pw(pma_checker_normal_entries_barrier_4_io_y_pw),
    .io_y_px(pma_checker_normal_entries_barrier_4_io_y_px),
    .io_y_pr(pma_checker_normal_entries_barrier_4_io_y_pr),
    .io_y_ppp(pma_checker_normal_entries_barrier_4_io_y_ppp),
    .io_y_pal(pma_checker_normal_entries_barrier_4_io_y_pal),
    .io_y_paa(pma_checker_normal_entries_barrier_4_io_y_paa),
    .io_y_eff(pma_checker_normal_entries_barrier_4_io_y_eff),
    .io_y_c(pma_checker_normal_entries_barrier_4_io_y_c)
  );
  OptimizationBarrier pma_checker_normal_entries_barrier_5 ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_normal_entries_barrier_5_io_x_ppn),
    .io_x_u(pma_checker_normal_entries_barrier_5_io_x_u),
    .io_x_ae(pma_checker_normal_entries_barrier_5_io_x_ae),
    .io_x_sw(pma_checker_normal_entries_barrier_5_io_x_sw),
    .io_x_sx(pma_checker_normal_entries_barrier_5_io_x_sx),
    .io_x_sr(pma_checker_normal_entries_barrier_5_io_x_sr),
    .io_x_pw(pma_checker_normal_entries_barrier_5_io_x_pw),
    .io_x_px(pma_checker_normal_entries_barrier_5_io_x_px),
    .io_x_pr(pma_checker_normal_entries_barrier_5_io_x_pr),
    .io_x_ppp(pma_checker_normal_entries_barrier_5_io_x_ppp),
    .io_x_pal(pma_checker_normal_entries_barrier_5_io_x_pal),
    .io_x_paa(pma_checker_normal_entries_barrier_5_io_x_paa),
    .io_x_eff(pma_checker_normal_entries_barrier_5_io_x_eff),
    .io_x_c(pma_checker_normal_entries_barrier_5_io_x_c),
    .io_y_ppn(pma_checker_normal_entries_barrier_5_io_y_ppn),
    .io_y_u(pma_checker_normal_entries_barrier_5_io_y_u),
    .io_y_ae(pma_checker_normal_entries_barrier_5_io_y_ae),
    .io_y_sw(pma_checker_normal_entries_barrier_5_io_y_sw),
    .io_y_sx(pma_checker_normal_entries_barrier_5_io_y_sx),
    .io_y_sr(pma_checker_normal_entries_barrier_5_io_y_sr),
    .io_y_pw(pma_checker_normal_entries_barrier_5_io_y_pw),
    .io_y_px(pma_checker_normal_entries_barrier_5_io_y_px),
    .io_y_pr(pma_checker_normal_entries_barrier_5_io_y_pr),
    .io_y_ppp(pma_checker_normal_entries_barrier_5_io_y_ppp),
    .io_y_pal(pma_checker_normal_entries_barrier_5_io_y_pal),
    .io_y_paa(pma_checker_normal_entries_barrier_5_io_y_paa),
    .io_y_eff(pma_checker_normal_entries_barrier_5_io_y_eff),
    .io_y_c(pma_checker_normal_entries_barrier_5_io_y_c)
  );
  OptimizationBarrier pma_checker_normal_entries_barrier_6 ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_normal_entries_barrier_6_io_x_ppn),
    .io_x_u(pma_checker_normal_entries_barrier_6_io_x_u),
    .io_x_ae(pma_checker_normal_entries_barrier_6_io_x_ae),
    .io_x_sw(pma_checker_normal_entries_barrier_6_io_x_sw),
    .io_x_sx(pma_checker_normal_entries_barrier_6_io_x_sx),
    .io_x_sr(pma_checker_normal_entries_barrier_6_io_x_sr),
    .io_x_pw(pma_checker_normal_entries_barrier_6_io_x_pw),
    .io_x_px(pma_checker_normal_entries_barrier_6_io_x_px),
    .io_x_pr(pma_checker_normal_entries_barrier_6_io_x_pr),
    .io_x_ppp(pma_checker_normal_entries_barrier_6_io_x_ppp),
    .io_x_pal(pma_checker_normal_entries_barrier_6_io_x_pal),
    .io_x_paa(pma_checker_normal_entries_barrier_6_io_x_paa),
    .io_x_eff(pma_checker_normal_entries_barrier_6_io_x_eff),
    .io_x_c(pma_checker_normal_entries_barrier_6_io_x_c),
    .io_y_ppn(pma_checker_normal_entries_barrier_6_io_y_ppn),
    .io_y_u(pma_checker_normal_entries_barrier_6_io_y_u),
    .io_y_ae(pma_checker_normal_entries_barrier_6_io_y_ae),
    .io_y_sw(pma_checker_normal_entries_barrier_6_io_y_sw),
    .io_y_sx(pma_checker_normal_entries_barrier_6_io_y_sx),
    .io_y_sr(pma_checker_normal_entries_barrier_6_io_y_sr),
    .io_y_pw(pma_checker_normal_entries_barrier_6_io_y_pw),
    .io_y_px(pma_checker_normal_entries_barrier_6_io_y_px),
    .io_y_pr(pma_checker_normal_entries_barrier_6_io_y_pr),
    .io_y_ppp(pma_checker_normal_entries_barrier_6_io_y_ppp),
    .io_y_pal(pma_checker_normal_entries_barrier_6_io_y_pal),
    .io_y_paa(pma_checker_normal_entries_barrier_6_io_y_paa),
    .io_y_eff(pma_checker_normal_entries_barrier_6_io_y_eff),
    .io_y_c(pma_checker_normal_entries_barrier_6_io_y_c)
  );
  OptimizationBarrier pma_checker_normal_entries_barrier_7 ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_normal_entries_barrier_7_io_x_ppn),
    .io_x_u(pma_checker_normal_entries_barrier_7_io_x_u),
    .io_x_ae(pma_checker_normal_entries_barrier_7_io_x_ae),
    .io_x_sw(pma_checker_normal_entries_barrier_7_io_x_sw),
    .io_x_sx(pma_checker_normal_entries_barrier_7_io_x_sx),
    .io_x_sr(pma_checker_normal_entries_barrier_7_io_x_sr),
    .io_x_pw(pma_checker_normal_entries_barrier_7_io_x_pw),
    .io_x_px(pma_checker_normal_entries_barrier_7_io_x_px),
    .io_x_pr(pma_checker_normal_entries_barrier_7_io_x_pr),
    .io_x_ppp(pma_checker_normal_entries_barrier_7_io_x_ppp),
    .io_x_pal(pma_checker_normal_entries_barrier_7_io_x_pal),
    .io_x_paa(pma_checker_normal_entries_barrier_7_io_x_paa),
    .io_x_eff(pma_checker_normal_entries_barrier_7_io_x_eff),
    .io_x_c(pma_checker_normal_entries_barrier_7_io_x_c),
    .io_y_ppn(pma_checker_normal_entries_barrier_7_io_y_ppn),
    .io_y_u(pma_checker_normal_entries_barrier_7_io_y_u),
    .io_y_ae(pma_checker_normal_entries_barrier_7_io_y_ae),
    .io_y_sw(pma_checker_normal_entries_barrier_7_io_y_sw),
    .io_y_sx(pma_checker_normal_entries_barrier_7_io_y_sx),
    .io_y_sr(pma_checker_normal_entries_barrier_7_io_y_sr),
    .io_y_pw(pma_checker_normal_entries_barrier_7_io_y_pw),
    .io_y_px(pma_checker_normal_entries_barrier_7_io_y_px),
    .io_y_pr(pma_checker_normal_entries_barrier_7_io_y_pr),
    .io_y_ppp(pma_checker_normal_entries_barrier_7_io_y_ppp),
    .io_y_pal(pma_checker_normal_entries_barrier_7_io_y_pal),
    .io_y_paa(pma_checker_normal_entries_barrier_7_io_y_paa),
    .io_y_eff(pma_checker_normal_entries_barrier_7_io_y_eff),
    .io_y_c(pma_checker_normal_entries_barrier_7_io_y_c)
  );
  OptimizationBarrier pma_checker_normal_entries_barrier_8 ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_normal_entries_barrier_8_io_x_ppn),
    .io_x_u(pma_checker_normal_entries_barrier_8_io_x_u),
    .io_x_ae(pma_checker_normal_entries_barrier_8_io_x_ae),
    .io_x_sw(pma_checker_normal_entries_barrier_8_io_x_sw),
    .io_x_sx(pma_checker_normal_entries_barrier_8_io_x_sx),
    .io_x_sr(pma_checker_normal_entries_barrier_8_io_x_sr),
    .io_x_pw(pma_checker_normal_entries_barrier_8_io_x_pw),
    .io_x_px(pma_checker_normal_entries_barrier_8_io_x_px),
    .io_x_pr(pma_checker_normal_entries_barrier_8_io_x_pr),
    .io_x_ppp(pma_checker_normal_entries_barrier_8_io_x_ppp),
    .io_x_pal(pma_checker_normal_entries_barrier_8_io_x_pal),
    .io_x_paa(pma_checker_normal_entries_barrier_8_io_x_paa),
    .io_x_eff(pma_checker_normal_entries_barrier_8_io_x_eff),
    .io_x_c(pma_checker_normal_entries_barrier_8_io_x_c),
    .io_y_ppn(pma_checker_normal_entries_barrier_8_io_y_ppn),
    .io_y_u(pma_checker_normal_entries_barrier_8_io_y_u),
    .io_y_ae(pma_checker_normal_entries_barrier_8_io_y_ae),
    .io_y_sw(pma_checker_normal_entries_barrier_8_io_y_sw),
    .io_y_sx(pma_checker_normal_entries_barrier_8_io_y_sx),
    .io_y_sr(pma_checker_normal_entries_barrier_8_io_y_sr),
    .io_y_pw(pma_checker_normal_entries_barrier_8_io_y_pw),
    .io_y_px(pma_checker_normal_entries_barrier_8_io_y_px),
    .io_y_pr(pma_checker_normal_entries_barrier_8_io_y_pr),
    .io_y_ppp(pma_checker_normal_entries_barrier_8_io_y_ppp),
    .io_y_pal(pma_checker_normal_entries_barrier_8_io_y_pal),
    .io_y_paa(pma_checker_normal_entries_barrier_8_io_y_paa),
    .io_y_eff(pma_checker_normal_entries_barrier_8_io_y_eff),
    .io_y_c(pma_checker_normal_entries_barrier_8_io_y_c)
  );
  OptimizationBarrier pma_checker_normal_entries_barrier_9 ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_normal_entries_barrier_9_io_x_ppn),
    .io_x_u(pma_checker_normal_entries_barrier_9_io_x_u),
    .io_x_ae(pma_checker_normal_entries_barrier_9_io_x_ae),
    .io_x_sw(pma_checker_normal_entries_barrier_9_io_x_sw),
    .io_x_sx(pma_checker_normal_entries_barrier_9_io_x_sx),
    .io_x_sr(pma_checker_normal_entries_barrier_9_io_x_sr),
    .io_x_pw(pma_checker_normal_entries_barrier_9_io_x_pw),
    .io_x_px(pma_checker_normal_entries_barrier_9_io_x_px),
    .io_x_pr(pma_checker_normal_entries_barrier_9_io_x_pr),
    .io_x_ppp(pma_checker_normal_entries_barrier_9_io_x_ppp),
    .io_x_pal(pma_checker_normal_entries_barrier_9_io_x_pal),
    .io_x_paa(pma_checker_normal_entries_barrier_9_io_x_paa),
    .io_x_eff(pma_checker_normal_entries_barrier_9_io_x_eff),
    .io_x_c(pma_checker_normal_entries_barrier_9_io_x_c),
    .io_y_ppn(pma_checker_normal_entries_barrier_9_io_y_ppn),
    .io_y_u(pma_checker_normal_entries_barrier_9_io_y_u),
    .io_y_ae(pma_checker_normal_entries_barrier_9_io_y_ae),
    .io_y_sw(pma_checker_normal_entries_barrier_9_io_y_sw),
    .io_y_sx(pma_checker_normal_entries_barrier_9_io_y_sx),
    .io_y_sr(pma_checker_normal_entries_barrier_9_io_y_sr),
    .io_y_pw(pma_checker_normal_entries_barrier_9_io_y_pw),
    .io_y_px(pma_checker_normal_entries_barrier_9_io_y_px),
    .io_y_pr(pma_checker_normal_entries_barrier_9_io_y_pr),
    .io_y_ppp(pma_checker_normal_entries_barrier_9_io_y_ppp),
    .io_y_pal(pma_checker_normal_entries_barrier_9_io_y_pal),
    .io_y_paa(pma_checker_normal_entries_barrier_9_io_y_paa),
    .io_y_eff(pma_checker_normal_entries_barrier_9_io_y_eff),
    .io_y_c(pma_checker_normal_entries_barrier_9_io_y_c)
  );
  OptimizationBarrier pma_checker_normal_entries_barrier_10 ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_normal_entries_barrier_10_io_x_ppn),
    .io_x_u(pma_checker_normal_entries_barrier_10_io_x_u),
    .io_x_ae(pma_checker_normal_entries_barrier_10_io_x_ae),
    .io_x_sw(pma_checker_normal_entries_barrier_10_io_x_sw),
    .io_x_sx(pma_checker_normal_entries_barrier_10_io_x_sx),
    .io_x_sr(pma_checker_normal_entries_barrier_10_io_x_sr),
    .io_x_pw(pma_checker_normal_entries_barrier_10_io_x_pw),
    .io_x_px(pma_checker_normal_entries_barrier_10_io_x_px),
    .io_x_pr(pma_checker_normal_entries_barrier_10_io_x_pr),
    .io_x_ppp(pma_checker_normal_entries_barrier_10_io_x_ppp),
    .io_x_pal(pma_checker_normal_entries_barrier_10_io_x_pal),
    .io_x_paa(pma_checker_normal_entries_barrier_10_io_x_paa),
    .io_x_eff(pma_checker_normal_entries_barrier_10_io_x_eff),
    .io_x_c(pma_checker_normal_entries_barrier_10_io_x_c),
    .io_y_ppn(pma_checker_normal_entries_barrier_10_io_y_ppn),
    .io_y_u(pma_checker_normal_entries_barrier_10_io_y_u),
    .io_y_ae(pma_checker_normal_entries_barrier_10_io_y_ae),
    .io_y_sw(pma_checker_normal_entries_barrier_10_io_y_sw),
    .io_y_sx(pma_checker_normal_entries_barrier_10_io_y_sx),
    .io_y_sr(pma_checker_normal_entries_barrier_10_io_y_sr),
    .io_y_pw(pma_checker_normal_entries_barrier_10_io_y_pw),
    .io_y_px(pma_checker_normal_entries_barrier_10_io_y_px),
    .io_y_pr(pma_checker_normal_entries_barrier_10_io_y_pr),
    .io_y_ppp(pma_checker_normal_entries_barrier_10_io_y_ppp),
    .io_y_pal(pma_checker_normal_entries_barrier_10_io_y_pal),
    .io_y_paa(pma_checker_normal_entries_barrier_10_io_y_paa),
    .io_y_eff(pma_checker_normal_entries_barrier_10_io_y_eff),
    .io_y_c(pma_checker_normal_entries_barrier_10_io_y_c)
  );
  OptimizationBarrier pma_checker_normal_entries_barrier_11 ( // @[package.scala 236:25]
    .io_x_ppn(pma_checker_normal_entries_barrier_11_io_x_ppn),
    .io_x_u(pma_checker_normal_entries_barrier_11_io_x_u),
    .io_x_ae(pma_checker_normal_entries_barrier_11_io_x_ae),
    .io_x_sw(pma_checker_normal_entries_barrier_11_io_x_sw),
    .io_x_sx(pma_checker_normal_entries_barrier_11_io_x_sx),
    .io_x_sr(pma_checker_normal_entries_barrier_11_io_x_sr),
    .io_x_pw(pma_checker_normal_entries_barrier_11_io_x_pw),
    .io_x_px(pma_checker_normal_entries_barrier_11_io_x_px),
    .io_x_pr(pma_checker_normal_entries_barrier_11_io_x_pr),
    .io_x_ppp(pma_checker_normal_entries_barrier_11_io_x_ppp),
    .io_x_pal(pma_checker_normal_entries_barrier_11_io_x_pal),
    .io_x_paa(pma_checker_normal_entries_barrier_11_io_x_paa),
    .io_x_eff(pma_checker_normal_entries_barrier_11_io_x_eff),
    .io_x_c(pma_checker_normal_entries_barrier_11_io_x_c),
    .io_y_ppn(pma_checker_normal_entries_barrier_11_io_y_ppn),
    .io_y_u(pma_checker_normal_entries_barrier_11_io_y_u),
    .io_y_ae(pma_checker_normal_entries_barrier_11_io_y_ae),
    .io_y_sw(pma_checker_normal_entries_barrier_11_io_y_sw),
    .io_y_sx(pma_checker_normal_entries_barrier_11_io_y_sx),
    .io_y_sr(pma_checker_normal_entries_barrier_11_io_y_sr),
    .io_y_pw(pma_checker_normal_entries_barrier_11_io_y_pw),
    .io_y_px(pma_checker_normal_entries_barrier_11_io_y_px),
    .io_y_pr(pma_checker_normal_entries_barrier_11_io_y_pr),
    .io_y_ppp(pma_checker_normal_entries_barrier_11_io_y_ppp),
    .io_y_pal(pma_checker_normal_entries_barrier_11_io_y_pal),
    .io_y_paa(pma_checker_normal_entries_barrier_11_io_y_paa),
    .io_y_eff(pma_checker_normal_entries_barrier_11_io_y_eff),
    .io_y_c(pma_checker_normal_entries_barrier_11_io_y_c)
  );
  MaxPeriodFibonacciLFSR lfsr_prng ( // @[PRNG.scala 82:22]
    .clock(lfsr_prng_clock),
    .reset(lfsr_prng_reset),
    .io_increment(lfsr_prng_io_increment),
    .io_out_0(lfsr_prng_io_out_0),
    .io_out_1(lfsr_prng_io_out_1),
    .io_out_2(lfsr_prng_io_out_2),
    .io_out_3(lfsr_prng_io_out_3),
    .io_out_4(lfsr_prng_io_out_4),
    .io_out_5(lfsr_prng_io_out_5),
    .io_out_6(lfsr_prng_io_out_6),
    .io_out_7(lfsr_prng_io_out_7),
    .io_out_8(lfsr_prng_io_out_8),
    .io_out_9(lfsr_prng_io_out_9),
    .io_out_10(lfsr_prng_io_out_10),
    .io_out_11(lfsr_prng_io_out_11),
    .io_out_12(lfsr_prng_io_out_12),
    .io_out_13(lfsr_prng_io_out_13),
    .io_out_14(lfsr_prng_io_out_14),
    .io_out_15(lfsr_prng_io_out_15)
  );
  tag_array tag_array ( // @[DescribedSRAM.scala 23:26]
    .RW0_addr(tag_array_RW0_addr),
    .RW0_en(tag_array_RW0_en),
    .RW0_clk(tag_array_RW0_clk),
    .RW0_wmode(tag_array_RW0_wmode),
    .RW0_wdata_0(tag_array_RW0_wdata_0),
    .RW0_wdata_1(tag_array_RW0_wdata_1),
    .RW0_wdata_2(tag_array_RW0_wdata_2),
    .RW0_wdata_3(tag_array_RW0_wdata_3),
    .RW0_rdata_0(tag_array_RW0_rdata_0),
    .RW0_rdata_1(tag_array_RW0_rdata_1),
    .RW0_rdata_2(tag_array_RW0_rdata_2),
    .RW0_rdata_3(tag_array_RW0_rdata_3),
    .RW0_wmask_0(tag_array_RW0_wmask_0),
    .RW0_wmask_1(tag_array_RW0_wmask_1),
    .RW0_wmask_2(tag_array_RW0_wmask_2),
    .RW0_wmask_3(tag_array_RW0_wmask_3)
  );
  DCacheDataArray data ( // @[DCache.scala 130:20]
    .clock(data_clock),
    .io_req_valid(data_io_req_valid),
    .io_req_bits_addr(data_io_req_bits_addr),
    .io_req_bits_write(data_io_req_bits_write),
    .io_req_bits_wdata(data_io_req_bits_wdata),
    .io_req_bits_eccMask(data_io_req_bits_eccMask),
    .io_req_bits_way_en(data_io_req_bits_way_en),
    .io_resp_0(data_io_resp_0),
    .io_resp_1(data_io_resp_1),
    .io_resp_2(data_io_resp_2),
    .io_resp_3(data_io_resp_3)
  );
  AMOALU amoalu ( // @[DCache.scala 881:26]
    .io_mask(amoalu_io_mask),
    .io_cmd(amoalu_io_cmd),
    .io_lhs(amoalu_io_lhs),
    .io_rhs(amoalu_io_rhs),
    .io_out(amoalu_io_out)
  );
  assign tlb_io_req_ready = tlb_state == 2'h0; // @[TLB.scala 337:25]
  assign tlb_io_resp_miss = tlb__io_resp_miss_T | tlb_multipleHits; // @[TLB.scala 350:41]
  assign tlb_io_resp_paddr = {tlb__ppn_T_53,tlb_mpu_physaddr_left}; // @[Cat.scala 29:58]
  assign tlb_io_resp_pf_ld = tlb__io_resp_pf_ld_T | tlb__io_resp_pf_ld_T_2; // @[TLB.scala 338:41]
  assign tlb_io_resp_pf_st = tlb__io_resp_pf_st_T | tlb__io_resp_pf_st_T_2; // @[TLB.scala 339:48]
  assign tlb_io_resp_ae_ld = |tlb__io_resp_ae_ld_T; // @[TLB.scala 341:41]
  assign tlb_io_resp_ae_st = |tlb__io_resp_ae_st_T; // @[TLB.scala 342:41]
  assign tlb_io_resp_ma_ld = |tlb__io_resp_ma_ld_T; // @[TLB.scala 344:41]
  assign tlb_io_resp_ma_st = |tlb__io_resp_ma_st_T; // @[TLB.scala 345:41]
  assign tlb_io_resp_cacheable = |tlb__io_resp_cacheable_T; // @[TLB.scala 347:41]
  assign tlb_io_ptw_req_valid = tlb_state == 2'h1; // @[TLB.scala 353:29]
  assign tlb_io_ptw_req_bits_bits_addr = tlb_r_refill_tag; // @[TLB.scala 355:29]
  assign tlb_mpu_ppn_data_barrier_io_x_ppn = tlb_special_entry_data_0[34:15]; // @[TLB.scala 86:77]
  assign tlb_mpu_ppn_data_barrier_io_x_u = tlb_special_entry_data_0[14]; // @[TLB.scala 86:77]
  assign tlb_mpu_ppn_data_barrier_io_x_ae = tlb_special_entry_data_0[12]; // @[TLB.scala 86:77]
  assign tlb_mpu_ppn_data_barrier_io_x_sw = tlb_special_entry_data_0[11]; // @[TLB.scala 86:77]
  assign tlb_mpu_ppn_data_barrier_io_x_sx = tlb_special_entry_data_0[10]; // @[TLB.scala 86:77]
  assign tlb_mpu_ppn_data_barrier_io_x_sr = tlb_special_entry_data_0[9]; // @[TLB.scala 86:77]
  assign tlb_mpu_ppn_data_barrier_io_x_pw = tlb_special_entry_data_0[8]; // @[TLB.scala 86:77]
  assign tlb_mpu_ppn_data_barrier_io_x_px = tlb_special_entry_data_0[7]; // @[TLB.scala 86:77]
  assign tlb_mpu_ppn_data_barrier_io_x_pr = tlb_special_entry_data_0[6]; // @[TLB.scala 86:77]
  assign tlb_mpu_ppn_data_barrier_io_x_ppp = tlb_special_entry_data_0[5]; // @[TLB.scala 86:77]
  assign tlb_mpu_ppn_data_barrier_io_x_pal = tlb_special_entry_data_0[4]; // @[TLB.scala 86:77]
  assign tlb_mpu_ppn_data_barrier_io_x_paa = tlb_special_entry_data_0[3]; // @[TLB.scala 86:77]
  assign tlb_mpu_ppn_data_barrier_io_x_eff = tlb_special_entry_data_0[2]; // @[TLB.scala 86:77]
  assign tlb_mpu_ppn_data_barrier_io_x_c = tlb_special_entry_data_0[1]; // @[TLB.scala 86:77]
  assign tlb_pmp_io_prv = tlb_mpu_priv[1:0]; // @[TLB.scala 194:14]
  assign tlb_pmp_io_pmp_0_cfg_l = tlb_io_ptw_pmp_0_cfg_l; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_0_cfg_a = tlb_io_ptw_pmp_0_cfg_a; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_0_cfg_x = tlb_io_ptw_pmp_0_cfg_x; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_0_cfg_w = tlb_io_ptw_pmp_0_cfg_w; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_0_cfg_r = tlb_io_ptw_pmp_0_cfg_r; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_0_addr = tlb_io_ptw_pmp_0_addr; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_0_mask = tlb_io_ptw_pmp_0_mask; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_1_cfg_l = tlb_io_ptw_pmp_1_cfg_l; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_1_cfg_a = tlb_io_ptw_pmp_1_cfg_a; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_1_cfg_x = tlb_io_ptw_pmp_1_cfg_x; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_1_cfg_w = tlb_io_ptw_pmp_1_cfg_w; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_1_cfg_r = tlb_io_ptw_pmp_1_cfg_r; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_1_addr = tlb_io_ptw_pmp_1_addr; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_1_mask = tlb_io_ptw_pmp_1_mask; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_2_cfg_l = tlb_io_ptw_pmp_2_cfg_l; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_2_cfg_a = tlb_io_ptw_pmp_2_cfg_a; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_2_cfg_x = tlb_io_ptw_pmp_2_cfg_x; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_2_cfg_w = tlb_io_ptw_pmp_2_cfg_w; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_2_cfg_r = tlb_io_ptw_pmp_2_cfg_r; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_2_addr = tlb_io_ptw_pmp_2_addr; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_2_mask = tlb_io_ptw_pmp_2_mask; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_3_cfg_l = tlb_io_ptw_pmp_3_cfg_l; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_3_cfg_a = tlb_io_ptw_pmp_3_cfg_a; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_3_cfg_x = tlb_io_ptw_pmp_3_cfg_x; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_3_cfg_w = tlb_io_ptw_pmp_3_cfg_w; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_3_cfg_r = tlb_io_ptw_pmp_3_cfg_r; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_3_addr = tlb_io_ptw_pmp_3_addr; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_3_mask = tlb_io_ptw_pmp_3_mask; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_4_cfg_l = tlb_io_ptw_pmp_4_cfg_l; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_4_cfg_a = tlb_io_ptw_pmp_4_cfg_a; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_4_cfg_x = tlb_io_ptw_pmp_4_cfg_x; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_4_cfg_w = tlb_io_ptw_pmp_4_cfg_w; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_4_cfg_r = tlb_io_ptw_pmp_4_cfg_r; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_4_addr = tlb_io_ptw_pmp_4_addr; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_4_mask = tlb_io_ptw_pmp_4_mask; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_5_cfg_l = tlb_io_ptw_pmp_5_cfg_l; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_5_cfg_a = tlb_io_ptw_pmp_5_cfg_a; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_5_cfg_x = tlb_io_ptw_pmp_5_cfg_x; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_5_cfg_w = tlb_io_ptw_pmp_5_cfg_w; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_5_cfg_r = tlb_io_ptw_pmp_5_cfg_r; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_5_addr = tlb_io_ptw_pmp_5_addr; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_5_mask = tlb_io_ptw_pmp_5_mask; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_6_cfg_l = tlb_io_ptw_pmp_6_cfg_l; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_6_cfg_a = tlb_io_ptw_pmp_6_cfg_a; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_6_cfg_x = tlb_io_ptw_pmp_6_cfg_x; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_6_cfg_w = tlb_io_ptw_pmp_6_cfg_w; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_6_cfg_r = tlb_io_ptw_pmp_6_cfg_r; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_6_addr = tlb_io_ptw_pmp_6_addr; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_6_mask = tlb_io_ptw_pmp_6_mask; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_7_cfg_l = tlb_io_ptw_pmp_7_cfg_l; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_7_cfg_a = tlb_io_ptw_pmp_7_cfg_a; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_7_cfg_x = tlb_io_ptw_pmp_7_cfg_x; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_7_cfg_w = tlb_io_ptw_pmp_7_cfg_w; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_7_cfg_r = tlb_io_ptw_pmp_7_cfg_r; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_7_addr = tlb_io_ptw_pmp_7_addr; // @[TLB.scala 193:14]
  assign tlb_pmp_io_pmp_7_mask = tlb_io_ptw_pmp_7_mask; // @[TLB.scala 193:14]
  assign tlb_pmp_io_addr = tlb_mpu_physaddr[31:0]; // @[TLB.scala 191:15]
  assign tlb_pmp_io_size = tlb_io_req_bits_size; // @[TLB.scala 192:15]
  assign tlb_ppn_data_barrier_io_x_ppn = tlb__GEN_35[34:15]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_io_x_u = tlb__GEN_35[14]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_io_x_ae = tlb__GEN_35[12]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_io_x_sw = tlb__GEN_35[11]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_io_x_sx = tlb__GEN_35[10]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_io_x_sr = tlb__GEN_35[9]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_io_x_pw = tlb__GEN_35[8]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_io_x_px = tlb__GEN_35[7]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_io_x_pr = tlb__GEN_35[6]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_io_x_ppp = tlb__GEN_35[5]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_io_x_pal = tlb__GEN_35[4]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_io_x_paa = tlb__GEN_35[3]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_io_x_eff = tlb__GEN_35[2]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_io_x_c = tlb__GEN_35[1]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_1_io_x_ppn = tlb__GEN_39[34:15]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_1_io_x_u = tlb__GEN_39[14]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_1_io_x_ae = tlb__GEN_39[12]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_1_io_x_sw = tlb__GEN_39[11]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_1_io_x_sx = tlb__GEN_39[10]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_1_io_x_sr = tlb__GEN_39[9]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_1_io_x_pw = tlb__GEN_39[8]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_1_io_x_px = tlb__GEN_39[7]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_1_io_x_pr = tlb__GEN_39[6]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_1_io_x_ppp = tlb__GEN_39[5]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_1_io_x_pal = tlb__GEN_39[4]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_1_io_x_paa = tlb__GEN_39[3]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_1_io_x_eff = tlb__GEN_39[2]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_1_io_x_c = tlb__GEN_39[1]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_2_io_x_ppn = tlb__GEN_43[34:15]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_2_io_x_u = tlb__GEN_43[14]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_2_io_x_ae = tlb__GEN_43[12]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_2_io_x_sw = tlb__GEN_43[11]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_2_io_x_sx = tlb__GEN_43[10]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_2_io_x_sr = tlb__GEN_43[9]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_2_io_x_pw = tlb__GEN_43[8]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_2_io_x_px = tlb__GEN_43[7]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_2_io_x_pr = tlb__GEN_43[6]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_2_io_x_ppp = tlb__GEN_43[5]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_2_io_x_pal = tlb__GEN_43[4]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_2_io_x_paa = tlb__GEN_43[3]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_2_io_x_eff = tlb__GEN_43[2]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_2_io_x_c = tlb__GEN_43[1]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_3_io_x_ppn = tlb__GEN_47[34:15]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_3_io_x_u = tlb__GEN_47[14]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_3_io_x_ae = tlb__GEN_47[12]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_3_io_x_sw = tlb__GEN_47[11]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_3_io_x_sx = tlb__GEN_47[10]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_3_io_x_sr = tlb__GEN_47[9]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_3_io_x_pw = tlb__GEN_47[8]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_3_io_x_px = tlb__GEN_47[7]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_3_io_x_pr = tlb__GEN_47[6]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_3_io_x_ppp = tlb__GEN_47[5]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_3_io_x_pal = tlb__GEN_47[4]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_3_io_x_paa = tlb__GEN_47[3]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_3_io_x_eff = tlb__GEN_47[2]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_3_io_x_c = tlb__GEN_47[1]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_4_io_x_ppn = tlb__GEN_51[34:15]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_4_io_x_u = tlb__GEN_51[14]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_4_io_x_ae = tlb__GEN_51[12]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_4_io_x_sw = tlb__GEN_51[11]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_4_io_x_sx = tlb__GEN_51[10]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_4_io_x_sr = tlb__GEN_51[9]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_4_io_x_pw = tlb__GEN_51[8]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_4_io_x_px = tlb__GEN_51[7]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_4_io_x_pr = tlb__GEN_51[6]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_4_io_x_ppp = tlb__GEN_51[5]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_4_io_x_pal = tlb__GEN_51[4]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_4_io_x_paa = tlb__GEN_51[3]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_4_io_x_eff = tlb__GEN_51[2]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_4_io_x_c = tlb__GEN_51[1]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_5_io_x_ppn = tlb__GEN_55[34:15]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_5_io_x_u = tlb__GEN_55[14]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_5_io_x_ae = tlb__GEN_55[12]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_5_io_x_sw = tlb__GEN_55[11]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_5_io_x_sx = tlb__GEN_55[10]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_5_io_x_sr = tlb__GEN_55[9]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_5_io_x_pw = tlb__GEN_55[8]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_5_io_x_px = tlb__GEN_55[7]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_5_io_x_pr = tlb__GEN_55[6]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_5_io_x_ppp = tlb__GEN_55[5]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_5_io_x_pal = tlb__GEN_55[4]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_5_io_x_paa = tlb__GEN_55[3]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_5_io_x_eff = tlb__GEN_55[2]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_5_io_x_c = tlb__GEN_55[1]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_6_io_x_ppn = tlb__GEN_59[34:15]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_6_io_x_u = tlb__GEN_59[14]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_6_io_x_ae = tlb__GEN_59[12]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_6_io_x_sw = tlb__GEN_59[11]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_6_io_x_sx = tlb__GEN_59[10]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_6_io_x_sr = tlb__GEN_59[9]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_6_io_x_pw = tlb__GEN_59[8]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_6_io_x_px = tlb__GEN_59[7]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_6_io_x_pr = tlb__GEN_59[6]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_6_io_x_ppp = tlb__GEN_59[5]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_6_io_x_pal = tlb__GEN_59[4]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_6_io_x_paa = tlb__GEN_59[3]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_6_io_x_eff = tlb__GEN_59[2]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_6_io_x_c = tlb__GEN_59[1]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_7_io_x_ppn = tlb__GEN_63[34:15]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_7_io_x_u = tlb__GEN_63[14]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_7_io_x_ae = tlb__GEN_63[12]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_7_io_x_sw = tlb__GEN_63[11]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_7_io_x_sx = tlb__GEN_63[10]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_7_io_x_sr = tlb__GEN_63[9]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_7_io_x_pw = tlb__GEN_63[8]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_7_io_x_px = tlb__GEN_63[7]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_7_io_x_pr = tlb__GEN_63[6]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_7_io_x_ppp = tlb__GEN_63[5]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_7_io_x_pal = tlb__GEN_63[4]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_7_io_x_paa = tlb__GEN_63[3]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_7_io_x_eff = tlb__GEN_63[2]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_7_io_x_c = tlb__GEN_63[1]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_8_io_x_ppn = tlb_superpage_entries_0_data_0[34:15]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_8_io_x_u = tlb_superpage_entries_0_data_0[14]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_8_io_x_ae = tlb_superpage_entries_0_data_0[12]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_8_io_x_sw = tlb_superpage_entries_0_data_0[11]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_8_io_x_sx = tlb_superpage_entries_0_data_0[10]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_8_io_x_sr = tlb_superpage_entries_0_data_0[9]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_8_io_x_pw = tlb_superpage_entries_0_data_0[8]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_8_io_x_px = tlb_superpage_entries_0_data_0[7]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_8_io_x_pr = tlb_superpage_entries_0_data_0[6]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_8_io_x_ppp = tlb_superpage_entries_0_data_0[5]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_8_io_x_pal = tlb_superpage_entries_0_data_0[4]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_8_io_x_paa = tlb_superpage_entries_0_data_0[3]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_8_io_x_eff = tlb_superpage_entries_0_data_0[2]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_8_io_x_c = tlb_superpage_entries_0_data_0[1]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_9_io_x_ppn = tlb_superpage_entries_1_data_0[34:15]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_9_io_x_u = tlb_superpage_entries_1_data_0[14]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_9_io_x_ae = tlb_superpage_entries_1_data_0[12]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_9_io_x_sw = tlb_superpage_entries_1_data_0[11]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_9_io_x_sx = tlb_superpage_entries_1_data_0[10]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_9_io_x_sr = tlb_superpage_entries_1_data_0[9]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_9_io_x_pw = tlb_superpage_entries_1_data_0[8]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_9_io_x_px = tlb_superpage_entries_1_data_0[7]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_9_io_x_pr = tlb_superpage_entries_1_data_0[6]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_9_io_x_ppp = tlb_superpage_entries_1_data_0[5]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_9_io_x_pal = tlb_superpage_entries_1_data_0[4]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_9_io_x_paa = tlb_superpage_entries_1_data_0[3]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_9_io_x_eff = tlb_superpage_entries_1_data_0[2]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_9_io_x_c = tlb_superpage_entries_1_data_0[1]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_10_io_x_ppn = tlb_superpage_entries_2_data_0[34:15]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_10_io_x_u = tlb_superpage_entries_2_data_0[14]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_10_io_x_ae = tlb_superpage_entries_2_data_0[12]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_10_io_x_sw = tlb_superpage_entries_2_data_0[11]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_10_io_x_sx = tlb_superpage_entries_2_data_0[10]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_10_io_x_sr = tlb_superpage_entries_2_data_0[9]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_10_io_x_pw = tlb_superpage_entries_2_data_0[8]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_10_io_x_px = tlb_superpage_entries_2_data_0[7]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_10_io_x_pr = tlb_superpage_entries_2_data_0[6]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_10_io_x_ppp = tlb_superpage_entries_2_data_0[5]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_10_io_x_pal = tlb_superpage_entries_2_data_0[4]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_10_io_x_paa = tlb_superpage_entries_2_data_0[3]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_10_io_x_eff = tlb_superpage_entries_2_data_0[2]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_10_io_x_c = tlb_superpage_entries_2_data_0[1]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_11_io_x_ppn = tlb_superpage_entries_3_data_0[34:15]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_11_io_x_u = tlb_superpage_entries_3_data_0[14]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_11_io_x_ae = tlb_superpage_entries_3_data_0[12]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_11_io_x_sw = tlb_superpage_entries_3_data_0[11]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_11_io_x_sx = tlb_superpage_entries_3_data_0[10]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_11_io_x_sr = tlb_superpage_entries_3_data_0[9]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_11_io_x_pw = tlb_superpage_entries_3_data_0[8]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_11_io_x_px = tlb_superpage_entries_3_data_0[7]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_11_io_x_pr = tlb_superpage_entries_3_data_0[6]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_11_io_x_ppp = tlb_superpage_entries_3_data_0[5]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_11_io_x_pal = tlb_superpage_entries_3_data_0[4]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_11_io_x_paa = tlb_superpage_entries_3_data_0[3]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_11_io_x_eff = tlb_superpage_entries_3_data_0[2]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_11_io_x_c = tlb_superpage_entries_3_data_0[1]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_12_io_x_ppn = tlb_special_entry_data_0[34:15]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_12_io_x_u = tlb_special_entry_data_0[14]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_12_io_x_ae = tlb_special_entry_data_0[12]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_12_io_x_sw = tlb_special_entry_data_0[11]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_12_io_x_sx = tlb_special_entry_data_0[10]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_12_io_x_sr = tlb_special_entry_data_0[9]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_12_io_x_pw = tlb_special_entry_data_0[8]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_12_io_x_px = tlb_special_entry_data_0[7]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_12_io_x_pr = tlb_special_entry_data_0[6]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_12_io_x_ppp = tlb_special_entry_data_0[5]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_12_io_x_pal = tlb_special_entry_data_0[4]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_12_io_x_paa = tlb_special_entry_data_0[3]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_12_io_x_eff = tlb_special_entry_data_0[2]; // @[TLB.scala 86:77]
  assign tlb_ppn_data_barrier_12_io_x_c = tlb_special_entry_data_0[1]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_io_x_ppn = tlb__GEN_35[34:15]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_io_x_u = tlb__GEN_35[14]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_io_x_ae = tlb__GEN_35[12]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_io_x_sw = tlb__GEN_35[11]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_io_x_sx = tlb__GEN_35[10]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_io_x_sr = tlb__GEN_35[9]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_io_x_pw = tlb__GEN_35[8]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_io_x_px = tlb__GEN_35[7]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_io_x_pr = tlb__GEN_35[6]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_io_x_ppp = tlb__GEN_35[5]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_io_x_pal = tlb__GEN_35[4]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_io_x_paa = tlb__GEN_35[3]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_io_x_eff = tlb__GEN_35[2]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_io_x_c = tlb__GEN_35[1]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_1_io_x_ppn = tlb__GEN_39[34:15]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_1_io_x_u = tlb__GEN_39[14]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_1_io_x_ae = tlb__GEN_39[12]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_1_io_x_sw = tlb__GEN_39[11]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_1_io_x_sx = tlb__GEN_39[10]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_1_io_x_sr = tlb__GEN_39[9]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_1_io_x_pw = tlb__GEN_39[8]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_1_io_x_px = tlb__GEN_39[7]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_1_io_x_pr = tlb__GEN_39[6]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_1_io_x_ppp = tlb__GEN_39[5]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_1_io_x_pal = tlb__GEN_39[4]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_1_io_x_paa = tlb__GEN_39[3]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_1_io_x_eff = tlb__GEN_39[2]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_1_io_x_c = tlb__GEN_39[1]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_2_io_x_ppn = tlb__GEN_43[34:15]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_2_io_x_u = tlb__GEN_43[14]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_2_io_x_ae = tlb__GEN_43[12]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_2_io_x_sw = tlb__GEN_43[11]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_2_io_x_sx = tlb__GEN_43[10]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_2_io_x_sr = tlb__GEN_43[9]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_2_io_x_pw = tlb__GEN_43[8]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_2_io_x_px = tlb__GEN_43[7]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_2_io_x_pr = tlb__GEN_43[6]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_2_io_x_ppp = tlb__GEN_43[5]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_2_io_x_pal = tlb__GEN_43[4]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_2_io_x_paa = tlb__GEN_43[3]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_2_io_x_eff = tlb__GEN_43[2]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_2_io_x_c = tlb__GEN_43[1]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_3_io_x_ppn = tlb__GEN_47[34:15]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_3_io_x_u = tlb__GEN_47[14]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_3_io_x_ae = tlb__GEN_47[12]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_3_io_x_sw = tlb__GEN_47[11]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_3_io_x_sx = tlb__GEN_47[10]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_3_io_x_sr = tlb__GEN_47[9]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_3_io_x_pw = tlb__GEN_47[8]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_3_io_x_px = tlb__GEN_47[7]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_3_io_x_pr = tlb__GEN_47[6]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_3_io_x_ppp = tlb__GEN_47[5]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_3_io_x_pal = tlb__GEN_47[4]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_3_io_x_paa = tlb__GEN_47[3]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_3_io_x_eff = tlb__GEN_47[2]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_3_io_x_c = tlb__GEN_47[1]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_4_io_x_ppn = tlb__GEN_51[34:15]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_4_io_x_u = tlb__GEN_51[14]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_4_io_x_ae = tlb__GEN_51[12]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_4_io_x_sw = tlb__GEN_51[11]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_4_io_x_sx = tlb__GEN_51[10]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_4_io_x_sr = tlb__GEN_51[9]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_4_io_x_pw = tlb__GEN_51[8]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_4_io_x_px = tlb__GEN_51[7]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_4_io_x_pr = tlb__GEN_51[6]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_4_io_x_ppp = tlb__GEN_51[5]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_4_io_x_pal = tlb__GEN_51[4]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_4_io_x_paa = tlb__GEN_51[3]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_4_io_x_eff = tlb__GEN_51[2]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_4_io_x_c = tlb__GEN_51[1]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_5_io_x_ppn = tlb__GEN_55[34:15]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_5_io_x_u = tlb__GEN_55[14]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_5_io_x_ae = tlb__GEN_55[12]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_5_io_x_sw = tlb__GEN_55[11]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_5_io_x_sx = tlb__GEN_55[10]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_5_io_x_sr = tlb__GEN_55[9]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_5_io_x_pw = tlb__GEN_55[8]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_5_io_x_px = tlb__GEN_55[7]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_5_io_x_pr = tlb__GEN_55[6]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_5_io_x_ppp = tlb__GEN_55[5]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_5_io_x_pal = tlb__GEN_55[4]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_5_io_x_paa = tlb__GEN_55[3]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_5_io_x_eff = tlb__GEN_55[2]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_5_io_x_c = tlb__GEN_55[1]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_6_io_x_ppn = tlb__GEN_59[34:15]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_6_io_x_u = tlb__GEN_59[14]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_6_io_x_ae = tlb__GEN_59[12]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_6_io_x_sw = tlb__GEN_59[11]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_6_io_x_sx = tlb__GEN_59[10]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_6_io_x_sr = tlb__GEN_59[9]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_6_io_x_pw = tlb__GEN_59[8]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_6_io_x_px = tlb__GEN_59[7]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_6_io_x_pr = tlb__GEN_59[6]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_6_io_x_ppp = tlb__GEN_59[5]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_6_io_x_pal = tlb__GEN_59[4]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_6_io_x_paa = tlb__GEN_59[3]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_6_io_x_eff = tlb__GEN_59[2]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_6_io_x_c = tlb__GEN_59[1]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_7_io_x_ppn = tlb__GEN_63[34:15]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_7_io_x_u = tlb__GEN_63[14]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_7_io_x_ae = tlb__GEN_63[12]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_7_io_x_sw = tlb__GEN_63[11]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_7_io_x_sx = tlb__GEN_63[10]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_7_io_x_sr = tlb__GEN_63[9]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_7_io_x_pw = tlb__GEN_63[8]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_7_io_x_px = tlb__GEN_63[7]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_7_io_x_pr = tlb__GEN_63[6]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_7_io_x_ppp = tlb__GEN_63[5]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_7_io_x_pal = tlb__GEN_63[4]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_7_io_x_paa = tlb__GEN_63[3]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_7_io_x_eff = tlb__GEN_63[2]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_7_io_x_c = tlb__GEN_63[1]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_8_io_x_ppn = tlb_superpage_entries_0_data_0[34:15]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_8_io_x_u = tlb_superpage_entries_0_data_0[14]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_8_io_x_ae = tlb_superpage_entries_0_data_0[12]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_8_io_x_sw = tlb_superpage_entries_0_data_0[11]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_8_io_x_sx = tlb_superpage_entries_0_data_0[10]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_8_io_x_sr = tlb_superpage_entries_0_data_0[9]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_8_io_x_pw = tlb_superpage_entries_0_data_0[8]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_8_io_x_px = tlb_superpage_entries_0_data_0[7]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_8_io_x_pr = tlb_superpage_entries_0_data_0[6]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_8_io_x_ppp = tlb_superpage_entries_0_data_0[5]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_8_io_x_pal = tlb_superpage_entries_0_data_0[4]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_8_io_x_paa = tlb_superpage_entries_0_data_0[3]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_8_io_x_eff = tlb_superpage_entries_0_data_0[2]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_8_io_x_c = tlb_superpage_entries_0_data_0[1]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_9_io_x_ppn = tlb_superpage_entries_1_data_0[34:15]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_9_io_x_u = tlb_superpage_entries_1_data_0[14]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_9_io_x_ae = tlb_superpage_entries_1_data_0[12]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_9_io_x_sw = tlb_superpage_entries_1_data_0[11]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_9_io_x_sx = tlb_superpage_entries_1_data_0[10]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_9_io_x_sr = tlb_superpage_entries_1_data_0[9]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_9_io_x_pw = tlb_superpage_entries_1_data_0[8]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_9_io_x_px = tlb_superpage_entries_1_data_0[7]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_9_io_x_pr = tlb_superpage_entries_1_data_0[6]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_9_io_x_ppp = tlb_superpage_entries_1_data_0[5]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_9_io_x_pal = tlb_superpage_entries_1_data_0[4]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_9_io_x_paa = tlb_superpage_entries_1_data_0[3]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_9_io_x_eff = tlb_superpage_entries_1_data_0[2]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_9_io_x_c = tlb_superpage_entries_1_data_0[1]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_10_io_x_ppn = tlb_superpage_entries_2_data_0[34:15]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_10_io_x_u = tlb_superpage_entries_2_data_0[14]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_10_io_x_ae = tlb_superpage_entries_2_data_0[12]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_10_io_x_sw = tlb_superpage_entries_2_data_0[11]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_10_io_x_sx = tlb_superpage_entries_2_data_0[10]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_10_io_x_sr = tlb_superpage_entries_2_data_0[9]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_10_io_x_pw = tlb_superpage_entries_2_data_0[8]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_10_io_x_px = tlb_superpage_entries_2_data_0[7]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_10_io_x_pr = tlb_superpage_entries_2_data_0[6]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_10_io_x_ppp = tlb_superpage_entries_2_data_0[5]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_10_io_x_pal = tlb_superpage_entries_2_data_0[4]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_10_io_x_paa = tlb_superpage_entries_2_data_0[3]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_10_io_x_eff = tlb_superpage_entries_2_data_0[2]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_10_io_x_c = tlb_superpage_entries_2_data_0[1]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_11_io_x_ppn = tlb_superpage_entries_3_data_0[34:15]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_11_io_x_u = tlb_superpage_entries_3_data_0[14]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_11_io_x_ae = tlb_superpage_entries_3_data_0[12]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_11_io_x_sw = tlb_superpage_entries_3_data_0[11]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_11_io_x_sx = tlb_superpage_entries_3_data_0[10]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_11_io_x_sr = tlb_superpage_entries_3_data_0[9]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_11_io_x_pw = tlb_superpage_entries_3_data_0[8]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_11_io_x_px = tlb_superpage_entries_3_data_0[7]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_11_io_x_pr = tlb_superpage_entries_3_data_0[6]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_11_io_x_ppp = tlb_superpage_entries_3_data_0[5]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_11_io_x_pal = tlb_superpage_entries_3_data_0[4]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_11_io_x_paa = tlb_superpage_entries_3_data_0[3]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_11_io_x_eff = tlb_superpage_entries_3_data_0[2]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_11_io_x_c = tlb_superpage_entries_3_data_0[1]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_12_io_x_ppn = tlb_special_entry_data_0[34:15]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_12_io_x_u = tlb_special_entry_data_0[14]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_12_io_x_ae = tlb_special_entry_data_0[12]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_12_io_x_sw = tlb_special_entry_data_0[11]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_12_io_x_sx = tlb_special_entry_data_0[10]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_12_io_x_sr = tlb_special_entry_data_0[9]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_12_io_x_pw = tlb_special_entry_data_0[8]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_12_io_x_px = tlb_special_entry_data_0[7]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_12_io_x_pr = tlb_special_entry_data_0[6]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_12_io_x_ppp = tlb_special_entry_data_0[5]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_12_io_x_pal = tlb_special_entry_data_0[4]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_12_io_x_paa = tlb_special_entry_data_0[3]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_12_io_x_eff = tlb_special_entry_data_0[2]; // @[TLB.scala 86:77]
  assign tlb_entries_barrier_12_io_x_c = tlb_special_entry_data_0[1]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_io_x_ppn = tlb__GEN_35[34:15]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_io_x_u = tlb__GEN_35[14]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_io_x_ae = tlb__GEN_35[12]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_io_x_sw = tlb__GEN_35[11]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_io_x_sx = tlb__GEN_35[10]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_io_x_sr = tlb__GEN_35[9]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_io_x_pw = tlb__GEN_35[8]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_io_x_px = tlb__GEN_35[7]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_io_x_pr = tlb__GEN_35[6]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_io_x_ppp = tlb__GEN_35[5]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_io_x_pal = tlb__GEN_35[4]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_io_x_paa = tlb__GEN_35[3]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_io_x_eff = tlb__GEN_35[2]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_io_x_c = tlb__GEN_35[1]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_1_io_x_ppn = tlb__GEN_39[34:15]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_1_io_x_u = tlb__GEN_39[14]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_1_io_x_ae = tlb__GEN_39[12]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_1_io_x_sw = tlb__GEN_39[11]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_1_io_x_sx = tlb__GEN_39[10]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_1_io_x_sr = tlb__GEN_39[9]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_1_io_x_pw = tlb__GEN_39[8]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_1_io_x_px = tlb__GEN_39[7]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_1_io_x_pr = tlb__GEN_39[6]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_1_io_x_ppp = tlb__GEN_39[5]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_1_io_x_pal = tlb__GEN_39[4]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_1_io_x_paa = tlb__GEN_39[3]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_1_io_x_eff = tlb__GEN_39[2]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_1_io_x_c = tlb__GEN_39[1]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_2_io_x_ppn = tlb__GEN_43[34:15]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_2_io_x_u = tlb__GEN_43[14]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_2_io_x_ae = tlb__GEN_43[12]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_2_io_x_sw = tlb__GEN_43[11]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_2_io_x_sx = tlb__GEN_43[10]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_2_io_x_sr = tlb__GEN_43[9]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_2_io_x_pw = tlb__GEN_43[8]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_2_io_x_px = tlb__GEN_43[7]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_2_io_x_pr = tlb__GEN_43[6]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_2_io_x_ppp = tlb__GEN_43[5]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_2_io_x_pal = tlb__GEN_43[4]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_2_io_x_paa = tlb__GEN_43[3]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_2_io_x_eff = tlb__GEN_43[2]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_2_io_x_c = tlb__GEN_43[1]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_3_io_x_ppn = tlb__GEN_47[34:15]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_3_io_x_u = tlb__GEN_47[14]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_3_io_x_ae = tlb__GEN_47[12]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_3_io_x_sw = tlb__GEN_47[11]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_3_io_x_sx = tlb__GEN_47[10]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_3_io_x_sr = tlb__GEN_47[9]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_3_io_x_pw = tlb__GEN_47[8]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_3_io_x_px = tlb__GEN_47[7]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_3_io_x_pr = tlb__GEN_47[6]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_3_io_x_ppp = tlb__GEN_47[5]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_3_io_x_pal = tlb__GEN_47[4]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_3_io_x_paa = tlb__GEN_47[3]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_3_io_x_eff = tlb__GEN_47[2]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_3_io_x_c = tlb__GEN_47[1]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_4_io_x_ppn = tlb__GEN_51[34:15]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_4_io_x_u = tlb__GEN_51[14]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_4_io_x_ae = tlb__GEN_51[12]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_4_io_x_sw = tlb__GEN_51[11]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_4_io_x_sx = tlb__GEN_51[10]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_4_io_x_sr = tlb__GEN_51[9]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_4_io_x_pw = tlb__GEN_51[8]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_4_io_x_px = tlb__GEN_51[7]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_4_io_x_pr = tlb__GEN_51[6]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_4_io_x_ppp = tlb__GEN_51[5]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_4_io_x_pal = tlb__GEN_51[4]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_4_io_x_paa = tlb__GEN_51[3]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_4_io_x_eff = tlb__GEN_51[2]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_4_io_x_c = tlb__GEN_51[1]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_5_io_x_ppn = tlb__GEN_55[34:15]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_5_io_x_u = tlb__GEN_55[14]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_5_io_x_ae = tlb__GEN_55[12]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_5_io_x_sw = tlb__GEN_55[11]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_5_io_x_sx = tlb__GEN_55[10]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_5_io_x_sr = tlb__GEN_55[9]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_5_io_x_pw = tlb__GEN_55[8]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_5_io_x_px = tlb__GEN_55[7]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_5_io_x_pr = tlb__GEN_55[6]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_5_io_x_ppp = tlb__GEN_55[5]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_5_io_x_pal = tlb__GEN_55[4]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_5_io_x_paa = tlb__GEN_55[3]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_5_io_x_eff = tlb__GEN_55[2]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_5_io_x_c = tlb__GEN_55[1]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_6_io_x_ppn = tlb__GEN_59[34:15]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_6_io_x_u = tlb__GEN_59[14]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_6_io_x_ae = tlb__GEN_59[12]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_6_io_x_sw = tlb__GEN_59[11]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_6_io_x_sx = tlb__GEN_59[10]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_6_io_x_sr = tlb__GEN_59[9]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_6_io_x_pw = tlb__GEN_59[8]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_6_io_x_px = tlb__GEN_59[7]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_6_io_x_pr = tlb__GEN_59[6]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_6_io_x_ppp = tlb__GEN_59[5]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_6_io_x_pal = tlb__GEN_59[4]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_6_io_x_paa = tlb__GEN_59[3]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_6_io_x_eff = tlb__GEN_59[2]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_6_io_x_c = tlb__GEN_59[1]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_7_io_x_ppn = tlb__GEN_63[34:15]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_7_io_x_u = tlb__GEN_63[14]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_7_io_x_ae = tlb__GEN_63[12]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_7_io_x_sw = tlb__GEN_63[11]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_7_io_x_sx = tlb__GEN_63[10]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_7_io_x_sr = tlb__GEN_63[9]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_7_io_x_pw = tlb__GEN_63[8]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_7_io_x_px = tlb__GEN_63[7]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_7_io_x_pr = tlb__GEN_63[6]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_7_io_x_ppp = tlb__GEN_63[5]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_7_io_x_pal = tlb__GEN_63[4]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_7_io_x_paa = tlb__GEN_63[3]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_7_io_x_eff = tlb__GEN_63[2]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_7_io_x_c = tlb__GEN_63[1]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_8_io_x_ppn = tlb_superpage_entries_0_data_0[34:15]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_8_io_x_u = tlb_superpage_entries_0_data_0[14]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_8_io_x_ae = tlb_superpage_entries_0_data_0[12]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_8_io_x_sw = tlb_superpage_entries_0_data_0[11]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_8_io_x_sx = tlb_superpage_entries_0_data_0[10]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_8_io_x_sr = tlb_superpage_entries_0_data_0[9]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_8_io_x_pw = tlb_superpage_entries_0_data_0[8]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_8_io_x_px = tlb_superpage_entries_0_data_0[7]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_8_io_x_pr = tlb_superpage_entries_0_data_0[6]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_8_io_x_ppp = tlb_superpage_entries_0_data_0[5]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_8_io_x_pal = tlb_superpage_entries_0_data_0[4]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_8_io_x_paa = tlb_superpage_entries_0_data_0[3]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_8_io_x_eff = tlb_superpage_entries_0_data_0[2]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_8_io_x_c = tlb_superpage_entries_0_data_0[1]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_9_io_x_ppn = tlb_superpage_entries_1_data_0[34:15]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_9_io_x_u = tlb_superpage_entries_1_data_0[14]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_9_io_x_ae = tlb_superpage_entries_1_data_0[12]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_9_io_x_sw = tlb_superpage_entries_1_data_0[11]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_9_io_x_sx = tlb_superpage_entries_1_data_0[10]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_9_io_x_sr = tlb_superpage_entries_1_data_0[9]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_9_io_x_pw = tlb_superpage_entries_1_data_0[8]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_9_io_x_px = tlb_superpage_entries_1_data_0[7]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_9_io_x_pr = tlb_superpage_entries_1_data_0[6]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_9_io_x_ppp = tlb_superpage_entries_1_data_0[5]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_9_io_x_pal = tlb_superpage_entries_1_data_0[4]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_9_io_x_paa = tlb_superpage_entries_1_data_0[3]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_9_io_x_eff = tlb_superpage_entries_1_data_0[2]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_9_io_x_c = tlb_superpage_entries_1_data_0[1]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_10_io_x_ppn = tlb_superpage_entries_2_data_0[34:15]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_10_io_x_u = tlb_superpage_entries_2_data_0[14]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_10_io_x_ae = tlb_superpage_entries_2_data_0[12]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_10_io_x_sw = tlb_superpage_entries_2_data_0[11]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_10_io_x_sx = tlb_superpage_entries_2_data_0[10]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_10_io_x_sr = tlb_superpage_entries_2_data_0[9]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_10_io_x_pw = tlb_superpage_entries_2_data_0[8]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_10_io_x_px = tlb_superpage_entries_2_data_0[7]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_10_io_x_pr = tlb_superpage_entries_2_data_0[6]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_10_io_x_ppp = tlb_superpage_entries_2_data_0[5]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_10_io_x_pal = tlb_superpage_entries_2_data_0[4]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_10_io_x_paa = tlb_superpage_entries_2_data_0[3]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_10_io_x_eff = tlb_superpage_entries_2_data_0[2]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_10_io_x_c = tlb_superpage_entries_2_data_0[1]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_11_io_x_ppn = tlb_superpage_entries_3_data_0[34:15]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_11_io_x_u = tlb_superpage_entries_3_data_0[14]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_11_io_x_ae = tlb_superpage_entries_3_data_0[12]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_11_io_x_sw = tlb_superpage_entries_3_data_0[11]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_11_io_x_sx = tlb_superpage_entries_3_data_0[10]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_11_io_x_sr = tlb_superpage_entries_3_data_0[9]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_11_io_x_pw = tlb_superpage_entries_3_data_0[8]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_11_io_x_px = tlb_superpage_entries_3_data_0[7]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_11_io_x_pr = tlb_superpage_entries_3_data_0[6]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_11_io_x_ppp = tlb_superpage_entries_3_data_0[5]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_11_io_x_pal = tlb_superpage_entries_3_data_0[4]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_11_io_x_paa = tlb_superpage_entries_3_data_0[3]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_11_io_x_eff = tlb_superpage_entries_3_data_0[2]; // @[TLB.scala 86:77]
  assign tlb_normal_entries_barrier_11_io_x_c = tlb_superpage_entries_3_data_0[1]; // @[TLB.scala 86:77]
  assign pma_checker_mpu_ppn_data_barrier_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_mpu_ppn_data_barrier_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_mpu_ppn_data_barrier_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_mpu_ppn_data_barrier_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_mpu_ppn_data_barrier_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_mpu_ppn_data_barrier_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_mpu_ppn_data_barrier_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_mpu_ppn_data_barrier_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_mpu_ppn_data_barrier_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_mpu_ppn_data_barrier_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_mpu_ppn_data_barrier_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_mpu_ppn_data_barrier_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_mpu_ppn_data_barrier_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_mpu_ppn_data_barrier_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_pmp_io_prv = 2'h1; // @[TLB.scala 194:14]
  assign pma_checker_pmp_io_pmp_0_cfg_l = 1'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_0_cfg_a = 2'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_0_cfg_x = 1'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_0_cfg_w = 1'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_0_cfg_r = 1'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_0_addr = 30'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_0_mask = 32'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_1_cfg_l = 1'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_1_cfg_a = 2'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_1_cfg_x = 1'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_1_cfg_w = 1'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_1_cfg_r = 1'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_1_addr = 30'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_1_mask = 32'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_2_cfg_l = 1'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_2_cfg_a = 2'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_2_cfg_x = 1'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_2_cfg_w = 1'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_2_cfg_r = 1'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_2_addr = 30'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_2_mask = 32'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_3_cfg_l = 1'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_3_cfg_a = 2'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_3_cfg_x = 1'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_3_cfg_w = 1'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_3_cfg_r = 1'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_3_addr = 30'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_3_mask = 32'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_4_cfg_l = 1'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_4_cfg_a = 2'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_4_cfg_x = 1'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_4_cfg_w = 1'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_4_cfg_r = 1'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_4_addr = 30'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_4_mask = 32'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_5_cfg_l = 1'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_5_cfg_a = 2'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_5_cfg_x = 1'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_5_cfg_w = 1'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_5_cfg_r = 1'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_5_addr = 30'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_5_mask = 32'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_6_cfg_l = 1'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_6_cfg_a = 2'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_6_cfg_x = 1'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_6_cfg_w = 1'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_6_cfg_r = 1'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_6_addr = 30'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_6_mask = 32'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_7_cfg_l = 1'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_7_cfg_a = 2'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_7_cfg_x = 1'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_7_cfg_w = 1'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_7_cfg_r = 1'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_7_addr = 30'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_pmp_7_mask = 32'h0; // @[TLB.scala 193:14]
  assign pma_checker_pmp_io_addr = 32'h0; // @[TLB.scala 191:15]
  assign pma_checker_pmp_io_size = pma_checker_io_req_bits_size; // @[TLB.scala 192:15]
  assign pma_checker_ppn_data_barrier_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_1_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_1_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_1_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_1_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_1_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_1_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_1_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_1_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_1_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_1_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_1_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_1_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_1_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_1_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_2_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_2_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_2_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_2_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_2_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_2_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_2_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_2_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_2_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_2_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_2_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_2_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_2_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_2_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_3_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_3_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_3_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_3_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_3_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_3_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_3_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_3_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_3_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_3_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_3_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_3_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_3_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_3_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_4_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_4_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_4_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_4_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_4_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_4_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_4_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_4_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_4_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_4_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_4_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_4_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_4_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_4_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_5_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_5_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_5_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_5_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_5_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_5_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_5_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_5_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_5_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_5_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_5_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_5_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_5_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_5_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_6_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_6_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_6_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_6_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_6_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_6_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_6_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_6_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_6_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_6_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_6_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_6_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_6_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_6_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_7_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_7_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_7_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_7_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_7_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_7_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_7_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_7_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_7_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_7_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_7_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_7_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_7_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_7_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_8_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_8_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_8_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_8_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_8_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_8_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_8_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_8_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_8_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_8_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_8_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_8_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_8_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_8_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_9_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_9_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_9_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_9_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_9_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_9_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_9_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_9_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_9_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_9_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_9_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_9_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_9_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_9_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_10_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_10_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_10_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_10_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_10_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_10_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_10_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_10_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_10_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_10_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_10_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_10_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_10_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_10_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_11_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_11_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_11_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_11_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_11_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_11_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_11_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_11_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_11_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_11_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_11_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_11_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_11_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_11_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_12_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_12_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_12_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_12_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_12_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_12_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_12_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_12_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_12_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_12_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_12_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_12_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_12_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_ppn_data_barrier_12_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_1_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_1_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_1_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_1_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_1_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_1_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_1_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_1_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_1_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_1_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_1_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_1_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_1_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_1_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_2_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_2_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_2_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_2_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_2_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_2_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_2_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_2_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_2_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_2_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_2_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_2_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_2_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_2_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_3_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_3_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_3_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_3_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_3_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_3_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_3_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_3_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_3_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_3_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_3_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_3_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_3_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_3_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_4_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_4_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_4_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_4_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_4_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_4_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_4_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_4_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_4_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_4_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_4_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_4_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_4_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_4_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_5_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_5_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_5_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_5_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_5_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_5_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_5_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_5_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_5_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_5_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_5_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_5_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_5_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_5_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_6_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_6_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_6_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_6_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_6_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_6_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_6_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_6_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_6_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_6_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_6_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_6_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_6_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_6_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_7_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_7_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_7_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_7_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_7_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_7_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_7_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_7_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_7_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_7_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_7_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_7_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_7_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_7_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_8_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_8_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_8_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_8_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_8_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_8_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_8_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_8_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_8_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_8_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_8_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_8_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_8_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_8_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_9_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_9_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_9_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_9_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_9_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_9_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_9_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_9_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_9_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_9_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_9_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_9_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_9_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_9_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_10_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_10_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_10_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_10_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_10_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_10_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_10_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_10_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_10_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_10_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_10_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_10_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_10_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_10_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_11_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_11_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_11_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_11_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_11_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_11_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_11_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_11_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_11_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_11_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_11_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_11_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_11_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_11_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_12_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_12_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_12_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_12_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_12_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_12_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_12_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_12_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_12_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_12_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_12_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_12_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_12_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_entries_barrier_12_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_1_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_1_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_1_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_1_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_1_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_1_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_1_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_1_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_1_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_1_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_1_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_1_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_1_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_1_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_2_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_2_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_2_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_2_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_2_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_2_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_2_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_2_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_2_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_2_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_2_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_2_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_2_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_2_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_3_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_3_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_3_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_3_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_3_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_3_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_3_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_3_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_3_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_3_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_3_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_3_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_3_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_3_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_4_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_4_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_4_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_4_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_4_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_4_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_4_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_4_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_4_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_4_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_4_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_4_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_4_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_4_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_5_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_5_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_5_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_5_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_5_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_5_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_5_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_5_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_5_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_5_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_5_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_5_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_5_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_5_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_6_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_6_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_6_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_6_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_6_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_6_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_6_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_6_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_6_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_6_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_6_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_6_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_6_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_6_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_7_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_7_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_7_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_7_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_7_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_7_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_7_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_7_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_7_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_7_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_7_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_7_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_7_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_7_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_8_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_8_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_8_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_8_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_8_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_8_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_8_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_8_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_8_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_8_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_8_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_8_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_8_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_8_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_9_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_9_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_9_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_9_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_9_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_9_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_9_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_9_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_9_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_9_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_9_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_9_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_9_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_9_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_10_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_10_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_10_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_10_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_10_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_10_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_10_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_10_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_10_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_10_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_10_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_10_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_10_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_10_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_11_io_x_ppn = 20'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_11_io_x_u = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_11_io_x_ae = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_11_io_x_sw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_11_io_x_sx = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_11_io_x_sr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_11_io_x_pw = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_11_io_x_px = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_11_io_x_pr = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_11_io_x_ppp = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_11_io_x_pal = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_11_io_x_paa = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_11_io_x_eff = 1'h0; // @[TLB.scala 86:77]
  assign pma_checker_normal_entries_barrier_11_io_x_c = 1'h0; // @[TLB.scala 86:77]
  assign metaArb_io_in_4_ready = ~metaArb__grant_T_2; // @[Arbiter.scala 31:78]
  assign metaArb_io_in_6_ready = ~metaArb__grant_T_3; // @[Arbiter.scala 31:78]
  assign metaArb_io_in_7_ready = ~metaArb__grant_T_5; // @[Arbiter.scala 31:78]
  assign metaArb_io_out_valid = metaArb__io_out_valid_T | metaArb_io_in_7_valid; // @[Arbiter.scala 135:31]
  assign metaArb_io_out_bits_write = metaArb_io_in_0_valid | metaArb__GEN_29; // @[Arbiter.scala 126:27 Arbiter.scala 128:19]
  assign metaArb_io_out_bits_addr = metaArb_io_in_0_valid ? metaArb_io_in_0_bits_addr : metaArb__GEN_28; // @[Arbiter.scala 126:27 Arbiter.scala 128:19]
  assign metaArb_io_out_bits_idx = metaArb_io_in_0_valid ? metaArb_io_in_0_bits_idx : metaArb__GEN_27; // @[Arbiter.scala 126:27 Arbiter.scala 128:19]
  assign metaArb_io_out_bits_way_en = metaArb_io_in_0_valid ? 4'hf : metaArb__GEN_26; // @[Arbiter.scala 126:27 Arbiter.scala 128:19]
  assign metaArb_io_out_bits_data = metaArb_io_in_0_valid ? metaArb_io_in_0_bits_data : metaArb__GEN_25; // @[Arbiter.scala 126:27 Arbiter.scala 128:19]
  assign dataArb_io_in_1_ready = ~dataArb_io_in_0_valid; // @[Arbiter.scala 31:78]
  assign dataArb_io_in_2_ready = ~dataArb__grant_T; // @[Arbiter.scala 31:78]
  assign dataArb_io_in_3_ready = ~dataArb__grant_T_1; // @[Arbiter.scala 31:78]
  assign dataArb_io_out_valid = dataArb__io_out_valid_T | dataArb_io_in_3_valid; // @[Arbiter.scala 135:31]
  assign dataArb_io_out_bits_addr = dataArb_io_in_0_valid ? dataArb_io_in_0_bits_addr : dataArb__GEN_13; // @[Arbiter.scala 126:27 Arbiter.scala 128:19]
  assign dataArb_io_out_bits_write = dataArb_io_in_0_valid ? dataArb_io_in_0_bits_write : dataArb__GEN_12; // @[Arbiter.scala 126:27 Arbiter.scala 128:19]
  assign dataArb_io_out_bits_wdata = dataArb_io_in_0_valid ? dataArb_io_in_0_bits_wdata : dataArb__GEN_11; // @[Arbiter.scala 126:27 Arbiter.scala 128:19]
  assign dataArb_io_out_bits_eccMask = dataArb_io_in_0_valid ? dataArb_io_in_0_bits_eccMask : 8'hff; // @[Arbiter.scala 126:27 Arbiter.scala 128:19]
  assign dataArb_io_out_bits_way_en = dataArb_io_in_0_valid ? dataArb_io_in_0_bits_way_en : dataArb__GEN_8; // @[Arbiter.scala 126:27 Arbiter.scala 128:19]
  assign auto_out_a_valid = s2_valid_uncached_pending | _tl_out_a_valid_T_6; // @[DCache.scala 550:67]
  assign auto_out_a_bits_opcode = _s2_valid_cached_miss_T ? 3'h6 : _tl_out_a_bits_T_8_opcode; // @[DCache.scala 552:23]
  assign auto_out_a_bits_param = _s2_valid_cached_miss_T ? tl_out_a_bits_a_param : _tl_out_a_bits_T_8_param; // @[DCache.scala 552:23]
  assign auto_out_a_bits_size = _s2_valid_cached_miss_T ? 4'h6 : _tl_out_a_bits_T_8_size; // @[DCache.scala 552:23]
  assign auto_out_a_bits_source = _s2_valid_cached_miss_T ? 1'h0 : _tl_out_a_bits_T_8_source; // @[DCache.scala 552:23]
  assign auto_out_a_bits_address = _s2_valid_cached_miss_T ? tl_out_a_bits_a_address : _tl_out_a_bits_T_8_address; // @[DCache.scala 552:23]
  assign auto_out_a_bits_mask = _s2_valid_cached_miss_T ? 8'hff : _tl_out_a_bits_T_8_mask; // @[DCache.scala 552:23]
  assign auto_out_a_bits_data = _s2_valid_cached_miss_T ? 64'h0 : _tl_out_a_bits_T_8_data; // @[DCache.scala 552:23]
  assign auto_out_b_ready = metaArb_io_in_6_ready & (~(((block_probe_for_core_progress | block_probe_for_ordering) |
    s1_valid) | s2_valid)); // @[DCache.scala 713:44]
  assign auto_out_c_valid = _T_271 | _GEN_301; // @[DCache.scala 774:48 DCache.scala 775:22]
  assign auto_out_c_bits_opcode = _T_275 ? 3'h7 : _GEN_314; // @[DCache.scala 783:81 DCache.scala 784:21]
  assign auto_out_c_bits_param = _T_275 ? s2_shrink_param : _GEN_315; // @[DCache.scala 783:81 DCache.scala 784:21]
  assign auto_out_c_bits_size = _T_275 ? 4'h6 : probe_bits_size; // @[DCache.scala 783:81 DCache.scala 784:21]
  assign auto_out_c_bits_source = probe_bits_source; // @[Nodes.scala 1213:84 DCache.scala 797:26]
  assign auto_out_c_bits_address = probe_bits_address; // @[Nodes.scala 1213:84 DCache.scala 798:27]
  assign auto_out_c_bits_data = {s2_data_corrected_right,s2_data_corrected_left}; // @[Cat.scala 29:58]
  assign auto_out_d_ready = _T_259 ? 1'h0 : _GEN_232; // @[DCache.scala 695:68 DCache.scala 696:22]
  assign auto_out_e_valid = _T_257 ? 1'h0 : _tl_out_e_valid_T_2; // @[DCache.scala 665:51 DCache.scala 666:20 DCache.scala 657:18]
  assign auto_out_e_bits_sink = auto_out_d_bits_sink; // @[Nodes.scala 1213:84 LazyModule.scala 314:12]
  assign io_cpu_req_ready = _T_259 ? _GEN_233 : _GEN_31; // @[DCache.scala 695:68]
  assign io_cpu_s2_nack = ((s2_valid_no_xcpt & (~s2_dont_nack_uncached)) & (~s2_dont_nack_misc)) & (~
    s2_valid_hit_pre_data_ecc_and_waw); // @[DCache.scala 396:86]
  assign io_cpu_resp_valid = s2_valid_hit_pre_data_ecc_and_waw | doUncachedResp; // @[DCache.scala 848:51]
  assign io_cpu_resp_bits_addr = doUncachedResp ? s2_uncached_resp_addr : s2_req_addr; // @[DCache.scala 850:25 DCache.scala 853:27 DCache.scala 819:20]
  assign io_cpu_resp_bits_tag = s2_req_tag; // @[DCache.scala 819:20]
  assign io_cpu_resp_bits_cmd = s2_req_cmd; // @[DCache.scala 819:20]
  assign io_cpu_resp_bits_size = s2_req_size; // @[DCache.scala 819:20]
  assign io_cpu_resp_bits_signed = s2_req_signed; // @[DCache.scala 819:20]
  assign io_cpu_resp_bits_dprv = s2_req_dprv; // @[DCache.scala 819:20]
  assign io_cpu_resp_bits_data = _io_cpu_resp_bits_data_T_23 | _GEN_398; // @[DCache.scala 873:41]
  assign io_cpu_resp_bits_mask = 8'h0; // @[DCache.scala 819:20]
  assign io_cpu_resp_bits_replay = doUncachedResp; // @[DCache.scala 850:25 DCache.scala 852:29 DCache.scala 821:27]
  assign io_cpu_resp_bits_has_data = (((s2_req_cmd == 5'h0) | _c_cat_T_47) | _s2_write_T_3) | _s2_write_T_21; // @[Consts.scala 82:75]
  assign io_cpu_resp_bits_data_word_bypass = {io_cpu_resp_bits_data_right,io_cpu_resp_bits_data_shifted}; // @[Cat.scala 29:58]
  assign io_cpu_resp_bits_data_raw = {s2_data_corrected_right,s2_data_corrected_left}; // @[Cat.scala 29:58]
  assign io_cpu_resp_bits_store_data = pstore1_data; // @[DCache.scala 876:31]
  assign io_cpu_replay_next = _T_236 & grantIsUncachedData; // @[DCache.scala 849:41]
  assign io_cpu_s2_xcpt_ma_ld = io_cpu_s2_xcpt_REG & s2_tlb_xcpt_ma_ld; // @[DCache.scala 832:24]
  assign io_cpu_s2_xcpt_ma_st = io_cpu_s2_xcpt_REG & s2_tlb_xcpt_ma_st; // @[DCache.scala 832:24]
  assign io_cpu_s2_xcpt_pf_ld = io_cpu_s2_xcpt_REG & s2_tlb_xcpt_pf_ld; // @[DCache.scala 832:24]
  assign io_cpu_s2_xcpt_pf_st = io_cpu_s2_xcpt_REG & s2_tlb_xcpt_pf_st; // @[DCache.scala 832:24]
  assign io_cpu_s2_xcpt_ae_ld = io_cpu_s2_xcpt_REG & s2_tlb_xcpt_ae_ld; // @[DCache.scala 832:24]
  assign io_cpu_s2_xcpt_ae_st = io_cpu_s2_xcpt_REG & s2_tlb_xcpt_ae_st; // @[DCache.scala 832:24]
  assign io_cpu_ordered = ~(((s1_valid | s2_valid) | cached_grant_wait) | _s2_valid_cached_miss_T_2); // @[DCache.scala 829:21]
  assign io_cpu_perf_release = io_cpu_perf_release_last & _T_262; // @[Edges.scala 234:22]
  assign io_cpu_perf_grant = auto_out_d_valid & d_last; // @[DCache.scala 979:39]
  assign io_ptw_req_valid = tlb_io_ptw_req_valid; // @[DCache.scala 230:10]
  assign io_ptw_req_bits_bits_addr = tlb_io_ptw_req_bits_bits_addr; // @[DCache.scala 230:10]
  assign tlb_clock = gated_clock;
  assign tlb_reset = reset;
  assign tlb_io_req_valid = s1_valid_masked & s1_cmd_uses_tlb; // @[DCache.scala 232:71]
  assign tlb_io_req_bits_vaddr = s1_tlb_req_vaddr; // @[DCache.scala 233:19]
  assign tlb_io_req_bits_passthrough = s1_tlb_req_passthrough; // @[DCache.scala 233:19]
  assign tlb_io_req_bits_size = s1_tlb_req_size; // @[DCache.scala 233:19]
  assign tlb_io_req_bits_cmd = s1_tlb_req_cmd; // @[DCache.scala 233:19]
  assign tlb_io_sfence_valid = s1_valid_masked & s1_sfence; // @[DCache.scala 237:54]
  assign tlb_io_sfence_bits_rs1 = s1_req_size[0]; // @[DCache.scala 238:40]
  assign tlb_io_sfence_bits_rs2 = s1_req_size[1]; // @[DCache.scala 239:40]
  assign tlb_io_sfence_bits_addr = s1_req_addr[38:0]; // @[DCache.scala 241:27]
  assign tlb_io_ptw_req_ready = io_ptw_req_ready; // @[DCache.scala 230:10]
  assign tlb_io_ptw_resp_valid = io_ptw_resp_valid; // @[DCache.scala 230:10]
  assign tlb_io_ptw_resp_bits_ae = io_ptw_resp_bits_ae; // @[DCache.scala 230:10]
  assign tlb_io_ptw_resp_bits_pte_ppn = io_ptw_resp_bits_pte_ppn; // @[DCache.scala 230:10]
  assign tlb_io_ptw_resp_bits_pte_d = io_ptw_resp_bits_pte_d; // @[DCache.scala 230:10]
  assign tlb_io_ptw_resp_bits_pte_a = io_ptw_resp_bits_pte_a; // @[DCache.scala 230:10]
  assign tlb_io_ptw_resp_bits_pte_g = io_ptw_resp_bits_pte_g; // @[DCache.scala 230:10]
  assign tlb_io_ptw_resp_bits_pte_u = io_ptw_resp_bits_pte_u; // @[DCache.scala 230:10]
  assign tlb_io_ptw_resp_bits_pte_x = io_ptw_resp_bits_pte_x; // @[DCache.scala 230:10]
  assign tlb_io_ptw_resp_bits_pte_w = io_ptw_resp_bits_pte_w; // @[DCache.scala 230:10]
  assign tlb_io_ptw_resp_bits_pte_r = io_ptw_resp_bits_pte_r; // @[DCache.scala 230:10]
  assign tlb_io_ptw_resp_bits_pte_v = io_ptw_resp_bits_pte_v; // @[DCache.scala 230:10]
  assign tlb_io_ptw_resp_bits_level = io_ptw_resp_bits_level; // @[DCache.scala 230:10]
  assign tlb_io_ptw_resp_bits_homogeneous = io_ptw_resp_bits_homogeneous; // @[DCache.scala 230:10]
  assign tlb_io_ptw_ptbr_mode = io_ptw_ptbr_mode; // @[DCache.scala 230:10]
  assign tlb_io_ptw_status_debug = io_ptw_status_debug; // @[DCache.scala 230:10]
  assign tlb_io_ptw_status_dprv = io_ptw_status_dprv; // @[DCache.scala 230:10]
  assign tlb_io_ptw_status_mxr = io_ptw_status_mxr; // @[DCache.scala 230:10]
  assign tlb_io_ptw_status_sum = io_ptw_status_sum; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_0_cfg_l = io_ptw_pmp_0_cfg_l; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_0_cfg_a = io_ptw_pmp_0_cfg_a; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_0_cfg_x = io_ptw_pmp_0_cfg_x; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_0_cfg_w = io_ptw_pmp_0_cfg_w; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_0_cfg_r = io_ptw_pmp_0_cfg_r; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_0_addr = io_ptw_pmp_0_addr; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_0_mask = io_ptw_pmp_0_mask; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_1_cfg_l = io_ptw_pmp_1_cfg_l; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_1_cfg_a = io_ptw_pmp_1_cfg_a; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_1_cfg_x = io_ptw_pmp_1_cfg_x; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_1_cfg_w = io_ptw_pmp_1_cfg_w; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_1_cfg_r = io_ptw_pmp_1_cfg_r; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_1_addr = io_ptw_pmp_1_addr; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_1_mask = io_ptw_pmp_1_mask; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_2_cfg_l = io_ptw_pmp_2_cfg_l; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_2_cfg_a = io_ptw_pmp_2_cfg_a; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_2_cfg_x = io_ptw_pmp_2_cfg_x; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_2_cfg_w = io_ptw_pmp_2_cfg_w; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_2_cfg_r = io_ptw_pmp_2_cfg_r; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_2_addr = io_ptw_pmp_2_addr; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_2_mask = io_ptw_pmp_2_mask; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_3_cfg_l = io_ptw_pmp_3_cfg_l; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_3_cfg_a = io_ptw_pmp_3_cfg_a; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_3_cfg_x = io_ptw_pmp_3_cfg_x; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_3_cfg_w = io_ptw_pmp_3_cfg_w; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_3_cfg_r = io_ptw_pmp_3_cfg_r; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_3_addr = io_ptw_pmp_3_addr; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_3_mask = io_ptw_pmp_3_mask; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_4_cfg_l = io_ptw_pmp_4_cfg_l; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_4_cfg_a = io_ptw_pmp_4_cfg_a; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_4_cfg_x = io_ptw_pmp_4_cfg_x; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_4_cfg_w = io_ptw_pmp_4_cfg_w; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_4_cfg_r = io_ptw_pmp_4_cfg_r; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_4_addr = io_ptw_pmp_4_addr; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_4_mask = io_ptw_pmp_4_mask; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_5_cfg_l = io_ptw_pmp_5_cfg_l; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_5_cfg_a = io_ptw_pmp_5_cfg_a; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_5_cfg_x = io_ptw_pmp_5_cfg_x; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_5_cfg_w = io_ptw_pmp_5_cfg_w; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_5_cfg_r = io_ptw_pmp_5_cfg_r; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_5_addr = io_ptw_pmp_5_addr; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_5_mask = io_ptw_pmp_5_mask; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_6_cfg_l = io_ptw_pmp_6_cfg_l; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_6_cfg_a = io_ptw_pmp_6_cfg_a; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_6_cfg_x = io_ptw_pmp_6_cfg_x; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_6_cfg_w = io_ptw_pmp_6_cfg_w; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_6_cfg_r = io_ptw_pmp_6_cfg_r; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_6_addr = io_ptw_pmp_6_addr; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_6_mask = io_ptw_pmp_6_mask; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_7_cfg_l = io_ptw_pmp_7_cfg_l; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_7_cfg_a = io_ptw_pmp_7_cfg_a; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_7_cfg_x = io_ptw_pmp_7_cfg_x; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_7_cfg_w = io_ptw_pmp_7_cfg_w; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_7_cfg_r = io_ptw_pmp_7_cfg_r; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_7_addr = io_ptw_pmp_7_addr; // @[DCache.scala 230:10]
  assign tlb_io_ptw_pmp_7_mask = io_ptw_pmp_7_mask; // @[DCache.scala 230:10]
  assign pma_checker_io_req_bits_size = s1_req_size; // @[DCache.scala 248:27]
  assign lfsr_prng_clock = gated_clock;
  assign lfsr_prng_reset = reset;
  assign lfsr_prng_io_increment = _T_236 & _GEN_208; // @[DCache.scala 617:26 Replacement.scala 37:11]
  assign metaArb_io_in_0_valid = resetting; // @[DCache.scala 947:26]
  assign metaArb_io_in_0_bits_addr = metaArb_io_in_5_bits_addr; // @[DCache.scala 948:25]
  assign metaArb_io_in_0_bits_idx = metaArb_io_in_5_bits_idx; // @[DCache.scala 948:25]
  assign metaArb_io_in_0_bits_data = {2'h0,metaArb_io_in_2_bits_data_meta_tag}; // @[DCache.scala 951:103]
  assign metaArb_io_in_2_valid = s2_valid_hit_pre_data_ecc_and_waw & s2_update_meta; // @[DCache.scala 413:63]
  assign metaArb_io_in_2_bits_addr = {metaArb_io_in_1_bits_addr_right,metaArb_io_in_2_bits_addr_left}; // @[Cat.scala 29:58]
  assign metaArb_io_in_2_bits_idx = s2_vaddr[11:6]; // @[DCache.scala 416:40]
  assign metaArb_io_in_2_bits_way_en = s2_hit_valid ? s2_hit_way : _s2_victim_way_T_1; // @[DCache.scala 383:26]
  assign metaArb_io_in_2_bits_data = {s2_grow_param,metaArb_io_in_2_bits_data_meta_tag}; // @[DCache.scala 418:97]
  assign metaArb_io_in_3_valid = (grantIsCached & d_done) & (~auto_out_d_bits_denied); // @[DCache.scala 684:53]
  assign metaArb_io_in_3_bits_addr = {metaArb_io_in_1_bits_addr_right,metaArb_io_in_2_bits_addr_left}; // @[Cat.scala 29:58]
  assign metaArb_io_in_3_bits_idx = s2_vaddr[11:6]; // @[DCache.scala 687:40]
  assign metaArb_io_in_3_bits_way_en = s2_hit_valid ? s2_hit_way : _s2_victim_way_T_1; // @[DCache.scala 383:26]
  assign metaArb_io_in_3_bits_data = {metaArb_io_in_3_bits_data_meta_state,metaArb_io_in_2_bits_data_meta_tag}; // @[DCache.scala 689:134]
  assign metaArb_io_in_4_valid = _T_274 | _metaArb_io_in_4_valid_T_1; // @[package.scala 64:59]
  assign metaArb_io_in_4_bits_addr = {metaArb_io_in_1_bits_addr_right,metaArb_io_in_4_bits_addr_left}; // @[Cat.scala 29:58]
  assign metaArb_io_in_4_bits_idx = probe_bits_address[11:6]; // @[DCache.scala 1095:47]
  assign metaArb_io_in_4_bits_way_en = _T_275 ? s2_victim_way : s2_probe_way; // @[DCache.scala 783:81 DCache.scala 790:18 DCache.scala 735:14]
  assign metaArb_io_in_4_bits_data = {newCoh_state,metaArb_io_in_4_bits_data_meta_tag}; // @[DCache.scala 815:97]
  assign metaArb_io_in_5_bits_addr = {metaArb_io_in_1_bits_addr_right,metaArb_io_in_5_bits_addr_left}; // @[Cat.scala 29:58]
  assign metaArb_io_in_5_bits_idx = flushCounter[5:0]; // @[DCache.scala 918:44]
  assign metaArb_io_in_6_valid = _T_269 | _metaArb_io_in_6_valid_T_2; // @[DCache.scala 761:44 DCache.scala 762:30 DCache.scala 712:26]
  assign metaArb_io_in_6_bits_addr = _T_269 ? _metaArb_io_in_6_bits_addr_T_1 : _metaArb_io_in_6_bits_addr_T; // @[DCache.scala 761:44 DCache.scala 764:34 DCache.scala 716:30]
  assign metaArb_io_in_6_bits_idx = _T_269 ? probe_bits_address[11:6] : auto_out_b_bits_address[11:6]; // @[DCache.scala 761:44 DCache.scala 763:33 DCache.scala 715:29]
  assign metaArb_io_in_6_bits_way_en = metaArb_io_in_4_bits_way_en; // @[DCache.scala 717:32]
  assign metaArb_io_in_6_bits_data = metaArb_io_in_4_bits_data; // @[DCache.scala 718:30]
  assign metaArb_io_in_7_valid = io_cpu_req_valid; // @[DCache.scala 220:26]
  assign metaArb_io_in_7_bits_addr = io_cpu_req_bits_addr; // @[DCache.scala 223:30]
  assign metaArb_io_in_7_bits_idx = io_cpu_req_bits_addr[11:6]; // @[DCache.scala 222:52]
  assign metaArb_io_in_7_bits_way_en = metaArb_io_in_4_bits_way_en; // @[DCache.scala 224:32]
  assign metaArb_io_in_7_bits_data = metaArb_io_in_4_bits_data; // @[DCache.scala 225:30]
  assign tag_array_RW0_wdata_0 = metaArb_io_out_bits_data; // @[compatibility.scala 127:12 compatibility.scala 127:12]
  assign tag_array_RW0_wdata_1 = metaArb_io_out_bits_data; // @[compatibility.scala 127:12 compatibility.scala 127:12]
  assign tag_array_RW0_wdata_2 = metaArb_io_out_bits_data; // @[compatibility.scala 127:12 compatibility.scala 127:12]
  assign tag_array_RW0_wdata_3 = metaArb_io_out_bits_data; // @[compatibility.scala 127:12 compatibility.scala 127:12]
  assign tag_array_RW0_wmask_0 = metaArb_io_out_bits_way_en[0]; // @[DCache.scala 263:74]
  assign tag_array_RW0_wmask_1 = metaArb_io_out_bits_way_en[1]; // @[DCache.scala 263:74]
  assign tag_array_RW0_wmask_2 = metaArb_io_out_bits_way_en[2]; // @[DCache.scala 263:74]
  assign tag_array_RW0_wmask_3 = metaArb_io_out_bits_way_en[3]; // @[DCache.scala 263:74]
  assign data_clock = gated_clock;
  assign data_io_req_valid = dataArb_io_out_valid; // @[DCache.scala 133:15]
  assign data_io_req_bits_addr = dataArb_io_out_bits_addr; // @[DCache.scala 133:15]
  assign data_io_req_bits_write = dataArb_io_out_bits_write; // @[DCache.scala 133:15]
  assign data_io_req_bits_wdata = dataArb_io_out_bits_wdata; // @[DCache.scala 133:15]
  assign data_io_req_bits_eccMask = dataArb_io_out_bits_eccMask; // @[DCache.scala 133:15]
  assign data_io_req_bits_way_en = dataArb_io_out_bits_way_en; // @[DCache.scala 133:15]
  assign dataArb_io_in_0_valid = pstore_drain_structural | _pstore_drain_T_10; // @[DCache.scala 468:48]
  assign dataArb_io_in_0_bits_addr = _dataArb_io_in_0_bits_addr_T[11:0]; // @[DCache.scala 500:30]
  assign dataArb_io_in_0_bits_write = pstore_drain_structural | _pstore_drain_T_10; // @[DCache.scala 468:48]
  assign dataArb_io_in_0_bits_wdata = {dataArb_io_in_0_bits_wdata_right,dataArb_io_in_0_bits_wdata_left}; // @[Cat.scala 29:58]
  assign dataArb_io_in_0_bits_eccMask = {dataArb_io_in_0_bits_eccMask_right,dataArb_io_in_0_bits_eccMask_left}; // @[Cat.scala 29:58]
  assign dataArb_io_in_0_bits_way_en = pstore2_valid ? pstore2_way : pstore1_way; // @[DCache.scala 501:38]
  assign dataArb_io_in_1_valid = _T_259 ? _GEN_234 : _dataArb_io_in_1_valid_T_1; // @[DCache.scala 695:68 DCache.scala 664:26]
  assign dataArb_io_in_1_bits_addr = _dataArb_io_in_1_bits_addr_T_2[11:0]; // @[DCache.scala 671:32]
  assign dataArb_io_in_1_bits_write = _T_259 ? _GEN_235 : 1'h1; // @[DCache.scala 695:68 DCache.scala 670:33]
  assign dataArb_io_in_1_bits_wdata = {tl_d_data_encoded_right,tl_d_data_encoded_left}; // @[Cat.scala 29:58]
  assign dataArb_io_in_1_bits_way_en = s2_hit_valid ? s2_hit_way : _s2_victim_way_T_1; // @[DCache.scala 383:26]
  assign dataArb_io_in_2_valid = inWriteback & (releaseDataBeat < 10'h8); // @[DCache.scala 803:41]
  assign dataArb_io_in_2_bits_addr = _dataArb_io_in_2_bits_addr_T_1 | _GEN_397; // @[DCache.scala 806:72]
  assign dataArb_io_in_2_bits_wdata = dataArb_io_in_1_bits_wdata; // @[DCache.scala 804:25]
  assign dataArb_io_in_3_valid = io_cpu_req_valid & res; // @[DCache.scala 212:46]
  assign dataArb_io_in_3_bits_addr = io_cpu_req_bits_addr[11:0]; // @[DCache.scala 215:30]
  assign dataArb_io_in_3_bits_wdata = dataArb_io_in_1_bits_wdata; // @[DCache.scala 213:25]
  assign amoalu_io_mask = pstore1_mask; // @[DCache.scala 882:38]
  assign amoalu_io_cmd = pstore1_cmd; // @[DCache.scala 883:21]
  assign amoalu_io_lhs = {s2_data_corrected_right,s2_data_corrected_left}; // @[Cat.scala 29:58]
  assign amoalu_io_rhs = pstore1_data; // @[DCache.scala 885:37]
  assign tag_array_RW0_wmode = metaArb_io_out_bits_write;
  assign tag_array_RW0_clk = gated_clock;
  assign tag_array_RW0_en = s0_clk_en | _T_19;
  assign tag_array_RW0_addr = metaArb_io_out_bits_idx;
  always @(posedge tlb_clock) begin
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_7) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_0_tag <= tlb_r_refill_tag; // @[TLB.scala 118:14]
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_7) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_0_data_0 <= tlb__GEN_89;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_7) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_0_data_1 <= tlb__GEN_90;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_7) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_0_data_2 <= tlb__GEN_91;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_7) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_0_data_3 <= tlb__GEN_92;
          end
        end
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_sectored_entries_0_valid_0 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__T_59) begin // @[TLB.scala 135:68]
          tlb_sectored_entries_0_valid_0 <= tlb__GEN_673;
        end else begin
          tlb_sectored_entries_0_valid_0 <= tlb__GEN_669;
        end
      end else begin
        tlb_sectored_entries_0_valid_0 <= tlb__GEN_685;
      end
    end else if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        tlb_sectored_entries_0_valid_0 <= tlb__GEN_305;
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_sectored_entries_0_valid_1 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__T_59) begin // @[TLB.scala 135:68]
          tlb_sectored_entries_0_valid_1 <= tlb__GEN_674;
        end else begin
          tlb_sectored_entries_0_valid_1 <= tlb__GEN_670;
        end
      end else begin
        tlb_sectored_entries_0_valid_1 <= tlb__GEN_686;
      end
    end else if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        tlb_sectored_entries_0_valid_1 <= tlb__GEN_306;
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_sectored_entries_0_valid_2 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__T_59) begin // @[TLB.scala 135:68]
          tlb_sectored_entries_0_valid_2 <= tlb__GEN_675;
        end else begin
          tlb_sectored_entries_0_valid_2 <= tlb__GEN_671;
        end
      end else begin
        tlb_sectored_entries_0_valid_2 <= tlb__GEN_687;
      end
    end else if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        tlb_sectored_entries_0_valid_2 <= tlb__GEN_307;
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_sectored_entries_0_valid_3 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__T_59) begin // @[TLB.scala 135:68]
          tlb_sectored_entries_0_valid_3 <= tlb__GEN_676;
        end else begin
          tlb_sectored_entries_0_valid_3 <= tlb__GEN_672;
        end
      end else begin
        tlb_sectored_entries_0_valid_3 <= tlb__GEN_688;
      end
    end else if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        tlb_sectored_entries_0_valid_3 <= tlb__GEN_308;
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_9) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_1_tag <= tlb_r_refill_tag; // @[TLB.scala 118:14]
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_9) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_1_data_0 <= tlb__GEN_115;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_9) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_1_data_1 <= tlb__GEN_116;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_9) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_1_data_2 <= tlb__GEN_117;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_9) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_1_data_3 <= tlb__GEN_118;
          end
        end
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_sectored_entries_1_valid_0 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__T_198) begin // @[TLB.scala 135:68]
          tlb_sectored_entries_1_valid_0 <= tlb__GEN_701;
        end else begin
          tlb_sectored_entries_1_valid_0 <= tlb__GEN_697;
        end
      end else begin
        tlb_sectored_entries_1_valid_0 <= tlb__GEN_713;
      end
    end else if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        tlb_sectored_entries_1_valid_0 <= tlb__GEN_315;
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_sectored_entries_1_valid_1 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__T_198) begin // @[TLB.scala 135:68]
          tlb_sectored_entries_1_valid_1 <= tlb__GEN_702;
        end else begin
          tlb_sectored_entries_1_valid_1 <= tlb__GEN_698;
        end
      end else begin
        tlb_sectored_entries_1_valid_1 <= tlb__GEN_714;
      end
    end else if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        tlb_sectored_entries_1_valid_1 <= tlb__GEN_316;
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_sectored_entries_1_valid_2 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__T_198) begin // @[TLB.scala 135:68]
          tlb_sectored_entries_1_valid_2 <= tlb__GEN_703;
        end else begin
          tlb_sectored_entries_1_valid_2 <= tlb__GEN_699;
        end
      end else begin
        tlb_sectored_entries_1_valid_2 <= tlb__GEN_715;
      end
    end else if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        tlb_sectored_entries_1_valid_2 <= tlb__GEN_317;
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_sectored_entries_1_valid_3 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__T_198) begin // @[TLB.scala 135:68]
          tlb_sectored_entries_1_valid_3 <= tlb__GEN_704;
        end else begin
          tlb_sectored_entries_1_valid_3 <= tlb__GEN_700;
        end
      end else begin
        tlb_sectored_entries_1_valid_3 <= tlb__GEN_716;
      end
    end else if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        tlb_sectored_entries_1_valid_3 <= tlb__GEN_318;
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_11) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_2_tag <= tlb_r_refill_tag; // @[TLB.scala 118:14]
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_11) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_2_data_0 <= tlb__GEN_141;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_11) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_2_data_1 <= tlb__GEN_142;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_11) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_2_data_2 <= tlb__GEN_143;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_11) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_2_data_3 <= tlb__GEN_144;
          end
        end
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_sectored_entries_2_valid_0 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__T_337) begin // @[TLB.scala 135:68]
          tlb_sectored_entries_2_valid_0 <= tlb__GEN_729;
        end else begin
          tlb_sectored_entries_2_valid_0 <= tlb__GEN_725;
        end
      end else begin
        tlb_sectored_entries_2_valid_0 <= tlb__GEN_741;
      end
    end else if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        tlb_sectored_entries_2_valid_0 <= tlb__GEN_325;
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_sectored_entries_2_valid_1 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__T_337) begin // @[TLB.scala 135:68]
          tlb_sectored_entries_2_valid_1 <= tlb__GEN_730;
        end else begin
          tlb_sectored_entries_2_valid_1 <= tlb__GEN_726;
        end
      end else begin
        tlb_sectored_entries_2_valid_1 <= tlb__GEN_742;
      end
    end else if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        tlb_sectored_entries_2_valid_1 <= tlb__GEN_326;
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_sectored_entries_2_valid_2 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__T_337) begin // @[TLB.scala 135:68]
          tlb_sectored_entries_2_valid_2 <= tlb__GEN_731;
        end else begin
          tlb_sectored_entries_2_valid_2 <= tlb__GEN_727;
        end
      end else begin
        tlb_sectored_entries_2_valid_2 <= tlb__GEN_743;
      end
    end else if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        tlb_sectored_entries_2_valid_2 <= tlb__GEN_327;
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_sectored_entries_2_valid_3 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__T_337) begin // @[TLB.scala 135:68]
          tlb_sectored_entries_2_valid_3 <= tlb__GEN_732;
        end else begin
          tlb_sectored_entries_2_valid_3 <= tlb__GEN_728;
        end
      end else begin
        tlb_sectored_entries_2_valid_3 <= tlb__GEN_744;
      end
    end else if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        tlb_sectored_entries_2_valid_3 <= tlb__GEN_328;
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_13) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_3_tag <= tlb_r_refill_tag; // @[TLB.scala 118:14]
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_13) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_3_data_0 <= tlb__GEN_167;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_13) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_3_data_1 <= tlb__GEN_168;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_13) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_3_data_2 <= tlb__GEN_169;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_13) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_3_data_3 <= tlb__GEN_170;
          end
        end
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_sectored_entries_3_valid_0 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__T_476) begin // @[TLB.scala 135:68]
          tlb_sectored_entries_3_valid_0 <= tlb__GEN_757;
        end else begin
          tlb_sectored_entries_3_valid_0 <= tlb__GEN_753;
        end
      end else begin
        tlb_sectored_entries_3_valid_0 <= tlb__GEN_769;
      end
    end else if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        tlb_sectored_entries_3_valid_0 <= tlb__GEN_335;
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_sectored_entries_3_valid_1 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__T_476) begin // @[TLB.scala 135:68]
          tlb_sectored_entries_3_valid_1 <= tlb__GEN_758;
        end else begin
          tlb_sectored_entries_3_valid_1 <= tlb__GEN_754;
        end
      end else begin
        tlb_sectored_entries_3_valid_1 <= tlb__GEN_770;
      end
    end else if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        tlb_sectored_entries_3_valid_1 <= tlb__GEN_336;
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_sectored_entries_3_valid_2 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__T_476) begin // @[TLB.scala 135:68]
          tlb_sectored_entries_3_valid_2 <= tlb__GEN_759;
        end else begin
          tlb_sectored_entries_3_valid_2 <= tlb__GEN_755;
        end
      end else begin
        tlb_sectored_entries_3_valid_2 <= tlb__GEN_771;
      end
    end else if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        tlb_sectored_entries_3_valid_2 <= tlb__GEN_337;
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_sectored_entries_3_valid_3 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__T_476) begin // @[TLB.scala 135:68]
          tlb_sectored_entries_3_valid_3 <= tlb__GEN_760;
        end else begin
          tlb_sectored_entries_3_valid_3 <= tlb__GEN_756;
        end
      end else begin
        tlb_sectored_entries_3_valid_3 <= tlb__GEN_772;
      end
    end else if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        tlb_sectored_entries_3_valid_3 <= tlb__GEN_338;
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_15) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_4_tag <= tlb_r_refill_tag; // @[TLB.scala 118:14]
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_15) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_4_data_0 <= tlb__GEN_193;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_15) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_4_data_1 <= tlb__GEN_194;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_15) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_4_data_2 <= tlb__GEN_195;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_15) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_4_data_3 <= tlb__GEN_196;
          end
        end
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_sectored_entries_4_valid_0 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__T_615) begin // @[TLB.scala 135:68]
          tlb_sectored_entries_4_valid_0 <= tlb__GEN_785;
        end else begin
          tlb_sectored_entries_4_valid_0 <= tlb__GEN_781;
        end
      end else begin
        tlb_sectored_entries_4_valid_0 <= tlb__GEN_797;
      end
    end else if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        tlb_sectored_entries_4_valid_0 <= tlb__GEN_345;
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_sectored_entries_4_valid_1 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__T_615) begin // @[TLB.scala 135:68]
          tlb_sectored_entries_4_valid_1 <= tlb__GEN_786;
        end else begin
          tlb_sectored_entries_4_valid_1 <= tlb__GEN_782;
        end
      end else begin
        tlb_sectored_entries_4_valid_1 <= tlb__GEN_798;
      end
    end else if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        tlb_sectored_entries_4_valid_1 <= tlb__GEN_346;
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_sectored_entries_4_valid_2 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__T_615) begin // @[TLB.scala 135:68]
          tlb_sectored_entries_4_valid_2 <= tlb__GEN_787;
        end else begin
          tlb_sectored_entries_4_valid_2 <= tlb__GEN_783;
        end
      end else begin
        tlb_sectored_entries_4_valid_2 <= tlb__GEN_799;
      end
    end else if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        tlb_sectored_entries_4_valid_2 <= tlb__GEN_347;
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_sectored_entries_4_valid_3 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__T_615) begin // @[TLB.scala 135:68]
          tlb_sectored_entries_4_valid_3 <= tlb__GEN_788;
        end else begin
          tlb_sectored_entries_4_valid_3 <= tlb__GEN_784;
        end
      end else begin
        tlb_sectored_entries_4_valid_3 <= tlb__GEN_800;
      end
    end else if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        tlb_sectored_entries_4_valid_3 <= tlb__GEN_348;
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_17) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_5_tag <= tlb_r_refill_tag; // @[TLB.scala 118:14]
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_17) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_5_data_0 <= tlb__GEN_219;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_17) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_5_data_1 <= tlb__GEN_220;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_17) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_5_data_2 <= tlb__GEN_221;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_17) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_5_data_3 <= tlb__GEN_222;
          end
        end
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_sectored_entries_5_valid_0 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__T_754) begin // @[TLB.scala 135:68]
          tlb_sectored_entries_5_valid_0 <= tlb__GEN_813;
        end else begin
          tlb_sectored_entries_5_valid_0 <= tlb__GEN_809;
        end
      end else begin
        tlb_sectored_entries_5_valid_0 <= tlb__GEN_825;
      end
    end else if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        tlb_sectored_entries_5_valid_0 <= tlb__GEN_355;
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_sectored_entries_5_valid_1 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__T_754) begin // @[TLB.scala 135:68]
          tlb_sectored_entries_5_valid_1 <= tlb__GEN_814;
        end else begin
          tlb_sectored_entries_5_valid_1 <= tlb__GEN_810;
        end
      end else begin
        tlb_sectored_entries_5_valid_1 <= tlb__GEN_826;
      end
    end else if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        tlb_sectored_entries_5_valid_1 <= tlb__GEN_356;
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_sectored_entries_5_valid_2 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__T_754) begin // @[TLB.scala 135:68]
          tlb_sectored_entries_5_valid_2 <= tlb__GEN_815;
        end else begin
          tlb_sectored_entries_5_valid_2 <= tlb__GEN_811;
        end
      end else begin
        tlb_sectored_entries_5_valid_2 <= tlb__GEN_827;
      end
    end else if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        tlb_sectored_entries_5_valid_2 <= tlb__GEN_357;
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_sectored_entries_5_valid_3 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__T_754) begin // @[TLB.scala 135:68]
          tlb_sectored_entries_5_valid_3 <= tlb__GEN_816;
        end else begin
          tlb_sectored_entries_5_valid_3 <= tlb__GEN_812;
        end
      end else begin
        tlb_sectored_entries_5_valid_3 <= tlb__GEN_828;
      end
    end else if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        tlb_sectored_entries_5_valid_3 <= tlb__GEN_358;
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_19) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_6_tag <= tlb_r_refill_tag; // @[TLB.scala 118:14]
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_19) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_6_data_0 <= tlb__GEN_245;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_19) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_6_data_1 <= tlb__GEN_246;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_19) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_6_data_2 <= tlb__GEN_247;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_19) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_6_data_3 <= tlb__GEN_248;
          end
        end
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_sectored_entries_6_valid_0 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__T_893) begin // @[TLB.scala 135:68]
          tlb_sectored_entries_6_valid_0 <= tlb__GEN_841;
        end else begin
          tlb_sectored_entries_6_valid_0 <= tlb__GEN_837;
        end
      end else begin
        tlb_sectored_entries_6_valid_0 <= tlb__GEN_853;
      end
    end else if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        tlb_sectored_entries_6_valid_0 <= tlb__GEN_365;
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_sectored_entries_6_valid_1 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__T_893) begin // @[TLB.scala 135:68]
          tlb_sectored_entries_6_valid_1 <= tlb__GEN_842;
        end else begin
          tlb_sectored_entries_6_valid_1 <= tlb__GEN_838;
        end
      end else begin
        tlb_sectored_entries_6_valid_1 <= tlb__GEN_854;
      end
    end else if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        tlb_sectored_entries_6_valid_1 <= tlb__GEN_366;
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_sectored_entries_6_valid_2 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__T_893) begin // @[TLB.scala 135:68]
          tlb_sectored_entries_6_valid_2 <= tlb__GEN_843;
        end else begin
          tlb_sectored_entries_6_valid_2 <= tlb__GEN_839;
        end
      end else begin
        tlb_sectored_entries_6_valid_2 <= tlb__GEN_855;
      end
    end else if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        tlb_sectored_entries_6_valid_2 <= tlb__GEN_367;
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_sectored_entries_6_valid_3 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__T_893) begin // @[TLB.scala 135:68]
          tlb_sectored_entries_6_valid_3 <= tlb__GEN_844;
        end else begin
          tlb_sectored_entries_6_valid_3 <= tlb__GEN_840;
        end
      end else begin
        tlb_sectored_entries_6_valid_3 <= tlb__GEN_856;
      end
    end else if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        tlb_sectored_entries_6_valid_3 <= tlb__GEN_368;
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_21) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_7_tag <= tlb_r_refill_tag; // @[TLB.scala 118:14]
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_21) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_7_data_0 <= tlb__GEN_271;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_21) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_7_data_1 <= tlb__GEN_272;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_21) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_7_data_2 <= tlb__GEN_273;
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (!(tlb__T_2)) begin // @[TLB.scala 242:54]
          if (tlb__T_21) begin // @[TLB.scala 249:72]
            tlb_sectored_entries_7_data_3 <= tlb__GEN_274;
          end
        end
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_sectored_entries_7_valid_0 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__T_1032) begin // @[TLB.scala 135:68]
          tlb_sectored_entries_7_valid_0 <= tlb__GEN_869;
        end else begin
          tlb_sectored_entries_7_valid_0 <= tlb__GEN_865;
        end
      end else begin
        tlb_sectored_entries_7_valid_0 <= tlb__GEN_881;
      end
    end else if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        tlb_sectored_entries_7_valid_0 <= tlb__GEN_375;
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_sectored_entries_7_valid_1 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__T_1032) begin // @[TLB.scala 135:68]
          tlb_sectored_entries_7_valid_1 <= tlb__GEN_870;
        end else begin
          tlb_sectored_entries_7_valid_1 <= tlb__GEN_866;
        end
      end else begin
        tlb_sectored_entries_7_valid_1 <= tlb__GEN_882;
      end
    end else if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        tlb_sectored_entries_7_valid_1 <= tlb__GEN_376;
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_sectored_entries_7_valid_2 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__T_1032) begin // @[TLB.scala 135:68]
          tlb_sectored_entries_7_valid_2 <= tlb__GEN_871;
        end else begin
          tlb_sectored_entries_7_valid_2 <= tlb__GEN_867;
        end
      end else begin
        tlb_sectored_entries_7_valid_2 <= tlb__GEN_883;
      end
    end else if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        tlb_sectored_entries_7_valid_2 <= tlb__GEN_377;
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_sectored_entries_7_valid_3 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__T_1032) begin // @[TLB.scala 135:68]
          tlb_sectored_entries_7_valid_3 <= tlb__GEN_872;
        end else begin
          tlb_sectored_entries_7_valid_3 <= tlb__GEN_868;
        end
      end else begin
        tlb_sectored_entries_7_valid_3 <= tlb__GEN_884;
      end
    end else if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        tlb_sectored_entries_7_valid_3 <= tlb__GEN_378;
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (tlb__T_2) begin // @[TLB.scala 242:54]
          if (tlb__T_3) begin // @[TLB.scala 243:89]
            tlb_superpage_entries_0_level <= {{1'd0}, tlb__superpage_entries_0_level_T}; // @[TLB.scala 119:16]
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (tlb__T_2) begin // @[TLB.scala 242:54]
          if (tlb__T_3) begin // @[TLB.scala 243:89]
            tlb_superpage_entries_0_tag <= tlb_r_refill_tag; // @[TLB.scala 118:14]
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (tlb__T_2) begin // @[TLB.scala 242:54]
          if (tlb__T_3) begin // @[TLB.scala 243:89]
            tlb_superpage_entries_0_data_0 <= tlb__special_entry_data_0_T; // @[TLB.scala 123:15]
          end
        end
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_superpage_entries_0_valid_0 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__superpage_hits_T_9) begin // @[TLB.scala 129:23]
          tlb_superpage_entries_0_valid_0 <= 1'h0; // @[TLB.scala 126:38]
        end else begin
          tlb_superpage_entries_0_valid_0 <= tlb__GEN_491;
        end
      end else begin
        tlb_superpage_entries_0_valid_0 <= tlb__GEN_891;
      end
    end else begin
      tlb_superpage_entries_0_valid_0 <= tlb__GEN_491;
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (tlb__T_2) begin // @[TLB.scala 242:54]
          if (tlb__T_4) begin // @[TLB.scala 243:89]
            tlb_superpage_entries_1_level <= {{1'd0}, tlb__superpage_entries_0_level_T}; // @[TLB.scala 119:16]
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (tlb__T_2) begin // @[TLB.scala 242:54]
          if (tlb__T_4) begin // @[TLB.scala 243:89]
            tlb_superpage_entries_1_tag <= tlb_r_refill_tag; // @[TLB.scala 118:14]
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (tlb__T_2) begin // @[TLB.scala 242:54]
          if (tlb__T_4) begin // @[TLB.scala 243:89]
            tlb_superpage_entries_1_data_0 <= tlb__special_entry_data_0_T; // @[TLB.scala 123:15]
          end
        end
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_superpage_entries_1_valid_0 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__superpage_hits_T_23) begin // @[TLB.scala 129:23]
          tlb_superpage_entries_1_valid_0 <= 1'h0; // @[TLB.scala 126:38]
        end else begin
          tlb_superpage_entries_1_valid_0 <= tlb__GEN_495;
        end
      end else begin
        tlb_superpage_entries_1_valid_0 <= tlb__GEN_895;
      end
    end else begin
      tlb_superpage_entries_1_valid_0 <= tlb__GEN_495;
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (tlb__T_2) begin // @[TLB.scala 242:54]
          if (tlb__T_5) begin // @[TLB.scala 243:89]
            tlb_superpage_entries_2_level <= {{1'd0}, tlb__superpage_entries_0_level_T}; // @[TLB.scala 119:16]
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (tlb__T_2) begin // @[TLB.scala 242:54]
          if (tlb__T_5) begin // @[TLB.scala 243:89]
            tlb_superpage_entries_2_tag <= tlb_r_refill_tag; // @[TLB.scala 118:14]
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (tlb__T_2) begin // @[TLB.scala 242:54]
          if (tlb__T_5) begin // @[TLB.scala 243:89]
            tlb_superpage_entries_2_data_0 <= tlb__special_entry_data_0_T; // @[TLB.scala 123:15]
          end
        end
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_superpage_entries_2_valid_0 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__superpage_hits_T_37) begin // @[TLB.scala 129:23]
          tlb_superpage_entries_2_valid_0 <= 1'h0; // @[TLB.scala 126:38]
        end else begin
          tlb_superpage_entries_2_valid_0 <= tlb__GEN_499;
        end
      end else begin
        tlb_superpage_entries_2_valid_0 <= tlb__GEN_899;
      end
    end else begin
      tlb_superpage_entries_2_valid_0 <= tlb__GEN_499;
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (tlb__T_2) begin // @[TLB.scala 242:54]
          if (tlb__T_6) begin // @[TLB.scala 243:89]
            tlb_superpage_entries_3_level <= {{1'd0}, tlb__superpage_entries_0_level_T}; // @[TLB.scala 119:16]
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (tlb__T_2) begin // @[TLB.scala 242:54]
          if (tlb__T_6) begin // @[TLB.scala 243:89]
            tlb_superpage_entries_3_tag <= tlb_r_refill_tag; // @[TLB.scala 118:14]
          end
        end
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(tlb__T)) begin // @[TLB.scala 237:68]
        if (tlb__T_2) begin // @[TLB.scala 242:54]
          if (tlb__T_6) begin // @[TLB.scala 243:89]
            tlb_superpage_entries_3_data_0 <= tlb__special_entry_data_0_T; // @[TLB.scala 123:15]
          end
        end
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_superpage_entries_3_valid_0 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__superpage_hits_T_51) begin // @[TLB.scala 129:23]
          tlb_superpage_entries_3_valid_0 <= 1'h0; // @[TLB.scala 126:38]
        end else begin
          tlb_superpage_entries_3_valid_0 <= tlb__GEN_503;
        end
      end else begin
        tlb_superpage_entries_3_valid_0 <= tlb__GEN_903;
      end
    end else begin
      tlb_superpage_entries_3_valid_0 <= tlb__GEN_503;
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (tlb__T) begin // @[TLB.scala 237:68]
        tlb_special_entry_level <= tlb_io_ptw_resp_bits_level; // @[TLB.scala 119:16]
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (tlb__T) begin // @[TLB.scala 237:68]
        tlb_special_entry_tag <= tlb_r_refill_tag; // @[TLB.scala 118:14]
      end
    end
    if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (tlb__T) begin // @[TLB.scala 237:68]
        tlb_special_entry_data_0 <= tlb__special_entry_data_0_T; // @[TLB.scala 123:15]
      end
    end
    if (tlb__T_1326) begin // @[TLB.scala 388:34]
      tlb_special_entry_valid_0 <= 1'h0; // @[TLB.scala 126:38]
    end else if (tlb_io_sfence_valid) begin // @[TLB.scala 380:19]
      if (tlb_io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (tlb__hitsVec_T_106) begin // @[TLB.scala 129:23]
          tlb_special_entry_valid_0 <= 1'h0; // @[TLB.scala 126:38]
        end else begin
          tlb_special_entry_valid_0 <= tlb__GEN_487;
        end
      end else begin
        tlb_special_entry_valid_0 <= tlb__GEN_907;
      end
    end else begin
      tlb_special_entry_valid_0 <= tlb__GEN_487;
    end
    if (tlb_reset) begin // @[TLB.scala 169:18]
      tlb_state <= 2'h0; // @[TLB.scala 169:18]
    end else if (tlb_io_ptw_resp_valid) begin // @[TLB.scala 376:30]
      tlb_state <= 2'h0; // @[TLB.scala 377:13]
    end else if (tlb__T_45) begin // @[TLB.scala 373:39]
      tlb_state <= 2'h3; // @[TLB.scala 374:13]
    end else if (tlb__invalidate_refill_T) begin // @[TLB.scala 368:32]
      tlb_state <= tlb__GEN_660;
    end else begin
      tlb_state <= tlb__GEN_653;
    end
    if (tlb__T_42) begin // @[TLB.scala 359:38]
      tlb_r_refill_tag <= tlb_vpn; // @[TLB.scala 361:20]
    end
    if (tlb__T_42) begin // @[TLB.scala 359:38]
      if (tlb__r_superpage_repl_addr_T_3) begin // @[TLB.scala 407:8]
        tlb_r_superpage_repl_addr <= tlb__r_superpage_repl_addr_T_2;
      end else if (tlb__r_superpage_repl_addr_T_5) begin // @[Mux.scala 47:69]
        tlb_r_superpage_repl_addr <= 2'h0;
      end else if (tlb__r_superpage_repl_addr_T_6) begin // @[Mux.scala 47:69]
        tlb_r_superpage_repl_addr <= 2'h1;
      end else begin
        tlb_r_superpage_repl_addr <= tlb__r_superpage_repl_addr_T_9;
      end
    end
    if (tlb__T_42) begin // @[TLB.scala 359:38]
      if (tlb__r_sectored_repl_addr_T_7) begin // @[TLB.scala 407:8]
        tlb_r_sectored_repl_addr <= tlb__r_sectored_repl_addr_T_6;
      end else if (tlb__r_sectored_repl_addr_T_9) begin // @[Mux.scala 47:69]
        tlb_r_sectored_repl_addr <= 3'h0;
      end else if (tlb__r_sectored_repl_addr_T_10) begin // @[Mux.scala 47:69]
        tlb_r_sectored_repl_addr <= 3'h1;
      end else begin
        tlb_r_sectored_repl_addr <= tlb__r_sectored_repl_addr_T_21;
      end
    end
    if (tlb__T_42) begin // @[TLB.scala 359:38]
      tlb_r_sectored_hit_addr <= tlb__T_34; // @[TLB.scala 365:27]
    end
    if (tlb__T_42) begin // @[TLB.scala 359:38]
      tlb_r_sectored_hit <= tlb__T_30; // @[TLB.scala 366:22]
    end
    if (tlb__T_23) begin // @[TLB.scala 325:37]
      if (tlb__T_30) begin // @[TLB.scala 326:28]
        tlb_state_reg <= tlb__state_reg_T_16; // @[Replacement.scala 162:15]
      end
    end
    if (tlb__T_23) begin // @[TLB.scala 325:37]
      if (tlb__T_37) begin // @[TLB.scala 327:31]
        tlb_state_reg_1 <= tlb__state_reg_1_T_6; // @[Replacement.scala 162:15]
      end
    end
  end
  always @(posedge gated_clock) begin
    if (reset) begin // @[DCache.scala 159:21]
      s1_valid <= 1'h0; // @[DCache.scala 159:21]
    end else begin
      s1_valid <= s1_valid_x9; // @[DCache.scala 159:21]
    end
    if (reset) begin // @[DCache.scala 611:38]
      blockProbeAfterGrantCount <= 3'h0; // @[DCache.scala 611:38]
    end else if (_T_236) begin // @[DCache.scala 617:26]
      if (grantIsCached) begin // @[DCache.scala 618:26]
        if (d_last) begin // @[DCache.scala 621:20]
          blockProbeAfterGrantCount <= 3'h7; // @[DCache.scala 624:35]
        end else begin
          blockProbeAfterGrantCount <= _GEN_182;
        end
      end else begin
        blockProbeAfterGrantCount <= _GEN_182;
      end
    end else begin
      blockProbeAfterGrantCount <= _GEN_182;
    end
    if (reset) begin // @[DCache.scala 423:22]
      lrscCount <= 7'h0; // @[DCache.scala 423:22]
    end else if (s1_probe) begin // @[DCache.scala 435:19]
      lrscCount <= 7'h0; // @[DCache.scala 435:31]
    end else if (_T_215) begin // @[DCache.scala 434:43]
      lrscCount <= 7'h3; // @[DCache.scala 434:55]
    end else if (_lrscBackingOff_T) begin // @[DCache.scala 433:24]
      lrscCount <= _lrscCount_T_2; // @[DCache.scala 433:36]
    end else begin
      lrscCount <= _GEN_120;
    end
    if (reset) begin // @[DCache.scala 160:21]
      s1_probe <= 1'h0; // @[DCache.scala 160:21]
    end else if (_T_269) begin // @[DCache.scala 761:44]
      s1_probe <= _GEN_294;
    end else begin
      s1_probe <= s1_probe_x12; // @[DCache.scala 160:21]
    end
    if (reset) begin // @[DCache.scala 285:21]
      s2_probe <= 1'h0; // @[DCache.scala 285:21]
    end else begin
      s2_probe <= s1_probe; // @[DCache.scala 285:21]
    end
    if (reset) begin // @[DCache.scala 199:26]
      release_state <= 3'h0; // @[DCache.scala 199:26]
    end else if (_T_278) begin // @[DCache.scala 816:34]
      release_state <= 3'h0; // @[DCache.scala 816:50]
    end else if (_T_275) begin // @[DCache.scala 783:81]
      if (releaseDone) begin // @[DCache.scala 791:26]
        release_state <= 3'h6; // @[DCache.scala 791:42]
      end else begin
        release_state <= _GEN_321;
      end
    end else begin
      release_state <= _GEN_321;
    end
    if (reset) begin // @[DCache.scala 197:29]
      release_ack_wait <= 1'h0; // @[DCache.scala 197:29]
    end else if (_T_275) begin // @[DCache.scala 783:81]
      release_ack_wait <= _GEN_323;
    end else if (_T_236) begin // @[DCache.scala 617:26]
      if (!(grantIsCached)) begin // @[DCache.scala 618:26]
        release_ack_wait <= _GEN_204;
      end
    end
    if (_T_275) begin // @[DCache.scala 783:81]
      if (_T_277) begin // @[DCache.scala 792:41]
        release_ack_addr <= probe_bits_address; // @[DCache.scala 794:26]
      end
    end
    if (reset) begin // @[DCache.scala 610:28]
      grantInProgress <= 1'h0; // @[DCache.scala 610:28]
    end else if (_T_236) begin // @[DCache.scala 617:26]
      if (grantIsCached) begin // @[DCache.scala 618:26]
        if (d_last) begin // @[DCache.scala 621:20]
          grantInProgress <= 1'h0; // @[DCache.scala 623:25]
        end else begin
          grantInProgress <= 1'h1; // @[DCache.scala 619:23]
        end
      end
    end
    if (reset) begin // @[DCache.scala 283:21]
      s2_valid <= 1'h0; // @[DCache.scala 283:21]
    end else begin
      s2_valid <= s2_valid_x36; // @[DCache.scala 283:21]
    end
    if (s2_want_victimize) begin // @[DCache.scala 738:25]
      probe_bits_param <= 2'h0; // @[DCache.scala 742:18]
    end else if (s1_probe_x12) begin // @[Reg.scala 16:19]
      probe_bits_param <= auto_out_b_bits_param; // @[Reg.scala 16:23]
    end
    if (s2_want_victimize) begin // @[DCache.scala 738:25]
      probe_bits_size <= 4'h0; // @[DCache.scala 742:18]
    end else if (s1_probe_x12) begin // @[Reg.scala 16:19]
      probe_bits_size <= auto_out_b_bits_size; // @[Reg.scala 16:23]
    end
    if (s2_want_victimize) begin // @[DCache.scala 738:25]
      probe_bits_source <= 1'h0; // @[DCache.scala 742:18]
    end else if (s1_probe_x12) begin // @[Reg.scala 16:19]
      probe_bits_source <= auto_out_b_bits_source; // @[Reg.scala 16:23]
    end
    if (s2_want_victimize) begin // @[DCache.scala 738:25]
      probe_bits_address <= res_2_address; // @[DCache.scala 742:18]
    end else if (s1_probe_x12) begin // @[Reg.scala 16:19]
      probe_bits_address <= auto_out_b_bits_address; // @[Reg.scala 16:23]
    end
    if (s1_probe) begin // @[Reg.scala 16:19]
      s2_probe_state_state <= s1_meta_hit_state_state; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[Edges.scala 230:27]
      counter_1 <= 9'h0; // @[Edges.scala 230:27]
    end else if (_T_262) begin // @[Edges.scala 236:17]
      if (c_first) begin // @[Edges.scala 237:21]
        if (beats1_opdata_1) begin // @[Edges.scala 222:14]
          counter_1 <= beats1_decode_1;
        end else begin
          counter_1 <= 9'h0;
        end
      end else begin
        counter_1 <= counter1_1;
      end
    end
    s2_release_data_valid <= s1_release_data_valid & (~releaseRejected); // @[DCache.scala 724:64]
    if (s0_clk_en) begin // @[Reg.scala 16:19]
      s1_req_cmd <= io_cpu_req_bits_cmd; // @[Reg.scala 16:23]
    end
    if (_T_236) begin // @[DCache.scala 617:26]
      if (grantIsCached) begin // @[DCache.scala 618:26]
        s2_req_cmd <= _GEN_59;
      end else if (grantIsUncached) begin // @[DCache.scala 627:35]
        if (grantIsUncachedData) begin // @[DCache.scala 634:34]
          s2_req_cmd <= 5'h0; // @[DCache.scala 638:22]
        end else begin
          s2_req_cmd <= _GEN_59;
        end
      end else begin
        s2_req_cmd <= _GEN_59;
      end
    end else begin
      s2_req_cmd <= _GEN_59;
    end
    pstore1_held <= (pstore1_valid & pstore2_valid) & (~pstore_drain); // @[DCache.scala 472:88]
    if (_pstore1_cmd_T) begin // @[Reg.scala 16:19]
      pstore1_addr <= s1_req_addr; // @[Reg.scala 16:23]
    end
    if (s0_clk_en) begin // @[Reg.scala 16:19]
      s1_req_addr <= s0_req_addr; // @[Reg.scala 16:23]
    end
    if (_pstore1_cmd_T) begin // @[Reg.scala 16:19]
      if (_s1_write_T_1) begin // @[DCache.scala 279:20]
        pstore1_mask <= io_cpu_s1_data_mask;
      end else begin
        pstore1_mask <= s1_mask_xwr;
      end
    end
    if (s0_clk_en) begin // @[Reg.scala 16:19]
      s1_req_size <= io_cpu_req_bits_size; // @[Reg.scala 16:23]
    end
    pstore2_valid <= (pstore2_valid & _pstore1_held_T_9) | advance_pstore1; // @[DCache.scala 474:51]
    if (advance_pstore1) begin // @[Reg.scala 16:19]
      pstore2_addr <= pstore1_addr; // @[Reg.scala 16:23]
    end
    if (advance_pstore1) begin // @[DCache.scala 483:45]
      mask <= _pstore2_storegen_mask_mask_T_2; // @[DCache.scala 485:12]
    end
    s2_not_nacked_in_s1 <= ~s1_nack; // @[DCache.scala 287:37]
    if (s1_valid_not_nacked) begin // @[Reg.scala 16:19]
      s2_hit_state_state <= s1_meta_hit_state_state; // @[Reg.scala 16:23]
    end
    if (s0_clk_en) begin // @[Reg.scala 16:19]
      s1_req_tag <= io_cpu_req_bits_tag; // @[Reg.scala 16:23]
    end
    if (s0_clk_en) begin // @[Reg.scala 16:19]
      s1_req_signed <= io_cpu_req_bits_signed; // @[Reg.scala 16:23]
    end
    if (s0_clk_en) begin // @[Reg.scala 16:19]
      s1_req_dprv <= io_cpu_req_bits_dprv; // @[Reg.scala 16:23]
    end
    if (s0_clk_en) begin // @[Reg.scala 16:19]
      s1_tlb_req_vaddr <= s0_req_addr; // @[Reg.scala 16:23]
    end
    if (s0_clk_en) begin // @[Reg.scala 16:19]
      s1_tlb_req_passthrough <= s0_req_phys; // @[Reg.scala 16:23]
    end
    if (s0_clk_en) begin // @[Reg.scala 16:19]
      s1_tlb_req_size <= io_cpu_req_bits_size; // @[Reg.scala 16:23]
    end
    if (s0_clk_en) begin // @[Reg.scala 16:19]
      s1_tlb_req_cmd <= io_cpu_req_bits_cmd; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[DCache.scala 196:30]
      cached_grant_wait <= 1'h0; // @[DCache.scala 196:30]
    end else if (_T_236) begin // @[DCache.scala 617:26]
      if (grantIsCached) begin // @[DCache.scala 618:26]
        if (d_last) begin // @[DCache.scala 621:20]
          cached_grant_wait <= 1'h0; // @[DCache.scala 622:27]
        end else begin
          cached_grant_wait <= _GEN_180;
        end
      end else begin
        cached_grant_wait <= _GEN_180;
      end
    end else begin
      cached_grant_wait <= _GEN_180;
    end
    if (reset) begin // @[DCache.scala 206:33]
      uncachedInFlight_0 <= 1'h0; // @[DCache.scala 206:33]
    end else if (_T_236) begin // @[DCache.scala 617:26]
      if (grantIsCached) begin // @[DCache.scala 618:26]
        uncachedInFlight_0 <= _GEN_168;
      end else if (grantIsUncached) begin // @[DCache.scala 627:35]
        uncachedInFlight_0 <= _GEN_187;
      end else begin
        uncachedInFlight_0 <= _GEN_168;
      end
    end else begin
      uncachedInFlight_0 <= _GEN_168;
    end
    if (_T_228) begin // @[DCache.scala 575:26]
      if (s2_uncached) begin // @[DCache.scala 576:24]
        if (a_sel) begin // @[DCache.scala 578:18]
          uncachedReqs_0_addr <= s2_req_addr; // @[DCache.scala 580:13]
        end
      end
    end
    if (_T_228) begin // @[DCache.scala 575:26]
      if (s2_uncached) begin // @[DCache.scala 576:24]
        if (a_sel) begin // @[DCache.scala 578:18]
          uncachedReqs_0_tag <= s2_req_tag; // @[DCache.scala 580:13]
        end
      end
    end
    if (_T_228) begin // @[DCache.scala 575:26]
      if (s2_uncached) begin // @[DCache.scala 576:24]
        if (a_sel) begin // @[DCache.scala 578:18]
          uncachedReqs_0_size <= s2_req_size; // @[DCache.scala 580:13]
        end
      end
    end
    if (_T_228) begin // @[DCache.scala 575:26]
      if (s2_uncached) begin // @[DCache.scala 576:24]
        if (a_sel) begin // @[DCache.scala 578:18]
          uncachedReqs_0_signed <= s2_req_signed; // @[DCache.scala 580:13]
        end
      end
    end
    if (s0_clk_en) begin // @[Reg.scala 16:19]
      s1_did_read <= _s1_did_read_T_52; // @[Reg.scala 16:23]
    end
    if (s1_valid_not_nacked) begin // @[Reg.scala 16:19]
      s2_hit_way <= s1_meta_hit_way; // @[Reg.scala 16:23]
    end
    if (s1_valid_not_nacked) begin // @[Reg.scala 16:19]
      s2_victim_way_r <= s1_victim_way_x32; // @[Reg.scala 16:23]
    end
    if (s1_probe) begin // @[Reg.scala 16:19]
      s2_probe_way <= s1_meta_hit_way; // @[Reg.scala 16:23]
    end
    if (_T_236) begin // @[DCache.scala 617:26]
      if (grantIsCached) begin // @[DCache.scala 618:26]
        s2_req_addr <= _GEN_57;
      end else if (grantIsUncached) begin // @[DCache.scala 627:35]
        if (grantIsUncachedData) begin // @[DCache.scala 634:34]
          s2_req_addr <= {{8'd0}, _s2_req_addr_T_1}; // @[DCache.scala 642:23]
        end else begin
          s2_req_addr <= _GEN_57;
        end
      end else begin
        s2_req_addr <= _GEN_57;
      end
    end else begin
      s2_req_addr <= _GEN_57;
    end
    if (_T_236) begin // @[DCache.scala 617:26]
      if (grantIsCached) begin // @[DCache.scala 618:26]
        s2_req_tag <= _GEN_58;
      end else if (grantIsUncached) begin // @[DCache.scala 627:35]
        if (grantIsUncachedData) begin // @[DCache.scala 634:34]
          s2_req_tag <= uncachedReqs_0_tag; // @[DCache.scala 641:22]
        end else begin
          s2_req_tag <= _GEN_58;
        end
      end else begin
        s2_req_tag <= _GEN_58;
      end
    end else begin
      s2_req_tag <= _GEN_58;
    end
    if (_T_236) begin // @[DCache.scala 617:26]
      if (grantIsCached) begin // @[DCache.scala 618:26]
        s2_req_size <= _GEN_60;
      end else if (grantIsUncached) begin // @[DCache.scala 627:35]
        if (grantIsUncachedData) begin // @[DCache.scala 634:34]
          s2_req_size <= uncachedReqs_0_size; // @[DCache.scala 639:23]
        end else begin
          s2_req_size <= _GEN_60;
        end
      end else begin
        s2_req_size <= _GEN_60;
      end
    end else begin
      s2_req_size <= _GEN_60;
    end
    if (_T_236) begin // @[DCache.scala 617:26]
      if (grantIsCached) begin // @[DCache.scala 618:26]
        s2_req_signed <= _GEN_61;
      end else if (grantIsUncached) begin // @[DCache.scala 627:35]
        if (grantIsUncachedData) begin // @[DCache.scala 634:34]
          s2_req_signed <= uncachedReqs_0_signed; // @[DCache.scala 640:25]
        end else begin
          s2_req_signed <= _GEN_61;
        end
      end else begin
        s2_req_signed <= _GEN_61;
      end
    end else begin
      s2_req_signed <= _GEN_61;
    end
    if (s1_valid_not_nacked) begin // @[DCache.scala 297:48]
      s2_req_dprv <= s1_req_dprv; // @[DCache.scala 298:12]
    end
    if (s1_valid_not_nacked) begin // @[DCache.scala 297:48]
      s2_tlb_xcpt_pf_ld <= tlb_io_resp_pf_ld; // @[DCache.scala 300:17]
    end
    if (s1_valid_not_nacked) begin // @[DCache.scala 297:48]
      s2_tlb_xcpt_pf_st <= tlb_io_resp_pf_st; // @[DCache.scala 300:17]
    end
    if (s1_valid_not_nacked) begin // @[DCache.scala 297:48]
      s2_tlb_xcpt_ae_ld <= tlb_io_resp_ae_ld; // @[DCache.scala 300:17]
    end
    if (s1_valid_not_nacked) begin // @[DCache.scala 297:48]
      s2_tlb_xcpt_ae_st <= tlb_io_resp_ae_st; // @[DCache.scala 300:17]
    end
    if (s1_valid_not_nacked) begin // @[DCache.scala 297:48]
      s2_tlb_xcpt_ma_ld <= tlb_io_resp_ma_ld; // @[DCache.scala 300:17]
    end
    if (s1_valid_not_nacked) begin // @[DCache.scala 297:48]
      s2_tlb_xcpt_ma_st <= tlb_io_resp_ma_st; // @[DCache.scala 300:17]
    end
    if (s1_valid_not_nacked) begin // @[DCache.scala 297:48]
      s2_pma_cacheable <= tlb_io_resp_cacheable; // @[DCache.scala 301:12]
    end
    if (_T_236) begin // @[DCache.scala 617:26]
      if (!(grantIsCached)) begin // @[DCache.scala 618:26]
        if (grantIsUncached) begin // @[DCache.scala 627:35]
          if (grantIsUncachedData) begin // @[DCache.scala 634:34]
            s2_uncached_resp_addr <= uncachedReqs_0_addr; // @[DCache.scala 647:33]
          end
        end
      end
    end
    if (s1_valid_not_nacked) begin // @[Reg.scala 16:19]
      s2_vaddr_r <= s1_req_addr; // @[Reg.scala 16:23]
    end
    if (_T_259) begin // @[DCache.scala 695:68]
      if (auto_out_d_valid) begin // @[DCache.scala 698:29]
        blockUncachedGrant <= _T_256; // @[DCache.scala 702:28]
      end else begin
        blockUncachedGrant <= dataArb_io_out_valid; // @[DCache.scala 694:24]
      end
    end else begin
      blockUncachedGrant <= dataArb_io_out_valid; // @[DCache.scala 694:24]
    end
    if (reset) begin // @[Edges.scala 230:27]
      counter <= 9'h0; // @[Edges.scala 230:27]
    end else if (_T_236) begin // @[Edges.scala 236:17]
      if (d_first) begin // @[Edges.scala 237:21]
        if (beats1_opdata) begin // @[Edges.scala 222:14]
          counter <= beats1_decode;
        end else begin
          counter <= 9'h0;
        end
      end else begin
        counter <= counter1;
      end
    end
    if (en) begin // @[Reg.scala 16:19]
      s2_data <= _s2_data_T_15; // @[Reg.scala 16:23]
    end
    if (s1_valid_not_nacked) begin // @[Reg.scala 16:19]
      if (s1_victim_way_x32 == 2'h3) begin // @[package.scala 32:76]
        s2_victim_tag_r <= s1_meta_uncorrected_3_tag;
      end else if (s1_victim_way_x32 == 2'h2) begin // @[package.scala 32:76]
        s2_victim_tag_r <= s1_meta_uncorrected_2_tag;
      end else if (s1_victim_way_x32 == 2'h1) begin // @[package.scala 32:76]
        s2_victim_tag_r <= s1_meta_uncorrected_1_tag;
      end else begin
        s2_victim_tag_r <= s1_meta_uncorrected_0_tag;
      end
    end
    if (s1_valid_not_nacked) begin // @[Reg.scala 16:19]
      if (s1_victim_way_x32 == 2'h3) begin // @[package.scala 32:76]
        s2_victim_state_r_state <= s1_meta_uncorrected_3_coh_state;
      end else if (s1_victim_way_x32 == 2'h2) begin // @[package.scala 32:76]
        s2_victim_state_r_state <= s1_meta_uncorrected_2_coh_state;
      end else if (s1_victim_way_x32 == 2'h1) begin // @[package.scala 32:76]
        s2_victim_state_r_state <= s1_meta_uncorrected_1_coh_state;
      end else begin
        s2_victim_state_r_state <= s1_meta_uncorrected_0_coh_state;
      end
    end
    if (_T_211) begin // @[DCache.scala 429:99]
      lrscAddr <= s2_req_addr[39:6]; // @[DCache.scala 431:14]
    end
    if (_pstore1_cmd_T) begin // @[Reg.scala 16:19]
      pstore1_cmd <= s1_req_cmd; // @[Reg.scala 16:23]
    end
    if (_pstore1_cmd_T) begin // @[Reg.scala 16:19]
      pstore1_data <= io_cpu_s1_data_data; // @[Reg.scala 16:23]
    end
    if (_pstore1_cmd_T) begin // @[Reg.scala 16:19]
      pstore1_way <= s1_meta_hit_way; // @[Reg.scala 16:23]
    end
    if (_pstore1_cmd_T) begin // @[Reg.scala 16:19]
      pstore1_rmw_r <= _pstore1_rmw_T_50; // @[Reg.scala 16:23]
    end
    pstore_drain_on_miss_REG <= io_cpu_s2_nack; // @[DCache.scala 454:56]
    if (advance_pstore1) begin // @[Reg.scala 16:19]
      pstore2_way <= pstore1_way; // @[Reg.scala 16:23]
    end
    if (advance_pstore1) begin // @[Reg.scala 16:19]
      pstore2_storegen_data_left_left_left <= pstore1_storegen_data[7:0]; // @[Reg.scala 16:23]
    end
    if (advance_pstore1) begin // @[Reg.scala 16:19]
      pstore2_storegen_data_left_left_right <= pstore1_storegen_data[15:8]; // @[Reg.scala 16:23]
    end
    if (advance_pstore1) begin // @[Reg.scala 16:19]
      pstore2_storegen_data_left_right_left <= pstore1_storegen_data[23:16]; // @[Reg.scala 16:23]
    end
    if (advance_pstore1) begin // @[Reg.scala 16:19]
      pstore2_storegen_data_left_right_right <= pstore1_storegen_data[31:24]; // @[Reg.scala 16:23]
    end
    if (advance_pstore1) begin // @[Reg.scala 16:19]
      pstore2_storegen_data_right_left_left <= pstore1_storegen_data[39:32]; // @[Reg.scala 16:23]
    end
    if (advance_pstore1) begin // @[Reg.scala 16:19]
      pstore2_storegen_data_right_left_right <= pstore1_storegen_data[47:40]; // @[Reg.scala 16:23]
    end
    if (advance_pstore1) begin // @[Reg.scala 16:19]
      pstore2_storegen_data_right_right_left <= pstore1_storegen_data[55:48]; // @[Reg.scala 16:23]
    end
    if (advance_pstore1) begin // @[Reg.scala 16:19]
      pstore2_storegen_data_right_right_right <= pstore1_storegen_data[63:56]; // @[Reg.scala 16:23]
    end
    s1_release_data_valid <= dataArb_io_in_2_ready & dataArb_io_in_2_valid; // @[Decoupled.scala 40:37]
    io_cpu_s2_xcpt_REG <= tlb_io_req_valid & _s1_valid_not_nacked_T; // @[DCache.scala 831:65]
    doUncachedResp <= io_cpu_replay_next; // @[DCache.scala 847:27]
    if (reset) begin // @[DCache.scala 906:26]
      resetting <= 1'h0; // @[DCache.scala 906:26]
    end else if (resetting) begin // @[DCache.scala 952:20]
      if (flushDone) begin // @[DCache.scala 954:22]
        resetting <= 1'h0; // @[DCache.scala 955:17]
      end else begin
        resetting <= _GEN_341;
      end
    end else begin
      resetting <= _GEN_341;
    end
    REG <= reset; // @[compatibility.scala 260:56]
    if (reset) begin // @[DCache.scala 909:25]
      flushCounter <= 8'hc0; // @[DCache.scala 909:25]
    end else begin
      flushCounter <= _GEN_343[7:0];
    end
    if (reset) begin // @[Edges.scala 230:27]
      io_cpu_perf_release_counter <= 9'h0; // @[Edges.scala 230:27]
    end else if (_T_262) begin // @[Edges.scala 236:17]
      if (io_cpu_perf_release_first) begin // @[Edges.scala 237:21]
        if (beats1_opdata_1) begin // @[Edges.scala 222:14]
          io_cpu_perf_release_counter <= beats1_decode_1;
        end else begin
          io_cpu_perf_release_counter <= 9'h0;
        end
      end else begin
        io_cpu_perf_release_counter <= io_cpu_perf_release_counter1;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  tlb_sectored_entries_0_tag = _RAND_0[26:0];
  _RAND_1 = {2{`RANDOM}};
  tlb_sectored_entries_0_data_0 = _RAND_1[34:0];
  _RAND_2 = {2{`RANDOM}};
  tlb_sectored_entries_0_data_1 = _RAND_2[34:0];
  _RAND_3 = {2{`RANDOM}};
  tlb_sectored_entries_0_data_2 = _RAND_3[34:0];
  _RAND_4 = {2{`RANDOM}};
  tlb_sectored_entries_0_data_3 = _RAND_4[34:0];
  _RAND_5 = {1{`RANDOM}};
  tlb_sectored_entries_0_valid_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  tlb_sectored_entries_0_valid_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  tlb_sectored_entries_0_valid_2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  tlb_sectored_entries_0_valid_3 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  tlb_sectored_entries_1_tag = _RAND_9[26:0];
  _RAND_10 = {2{`RANDOM}};
  tlb_sectored_entries_1_data_0 = _RAND_10[34:0];
  _RAND_11 = {2{`RANDOM}};
  tlb_sectored_entries_1_data_1 = _RAND_11[34:0];
  _RAND_12 = {2{`RANDOM}};
  tlb_sectored_entries_1_data_2 = _RAND_12[34:0];
  _RAND_13 = {2{`RANDOM}};
  tlb_sectored_entries_1_data_3 = _RAND_13[34:0];
  _RAND_14 = {1{`RANDOM}};
  tlb_sectored_entries_1_valid_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  tlb_sectored_entries_1_valid_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  tlb_sectored_entries_1_valid_2 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  tlb_sectored_entries_1_valid_3 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  tlb_sectored_entries_2_tag = _RAND_18[26:0];
  _RAND_19 = {2{`RANDOM}};
  tlb_sectored_entries_2_data_0 = _RAND_19[34:0];
  _RAND_20 = {2{`RANDOM}};
  tlb_sectored_entries_2_data_1 = _RAND_20[34:0];
  _RAND_21 = {2{`RANDOM}};
  tlb_sectored_entries_2_data_2 = _RAND_21[34:0];
  _RAND_22 = {2{`RANDOM}};
  tlb_sectored_entries_2_data_3 = _RAND_22[34:0];
  _RAND_23 = {1{`RANDOM}};
  tlb_sectored_entries_2_valid_0 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  tlb_sectored_entries_2_valid_1 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  tlb_sectored_entries_2_valid_2 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  tlb_sectored_entries_2_valid_3 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  tlb_sectored_entries_3_tag = _RAND_27[26:0];
  _RAND_28 = {2{`RANDOM}};
  tlb_sectored_entries_3_data_0 = _RAND_28[34:0];
  _RAND_29 = {2{`RANDOM}};
  tlb_sectored_entries_3_data_1 = _RAND_29[34:0];
  _RAND_30 = {2{`RANDOM}};
  tlb_sectored_entries_3_data_2 = _RAND_30[34:0];
  _RAND_31 = {2{`RANDOM}};
  tlb_sectored_entries_3_data_3 = _RAND_31[34:0];
  _RAND_32 = {1{`RANDOM}};
  tlb_sectored_entries_3_valid_0 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  tlb_sectored_entries_3_valid_1 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  tlb_sectored_entries_3_valid_2 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  tlb_sectored_entries_3_valid_3 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  tlb_sectored_entries_4_tag = _RAND_36[26:0];
  _RAND_37 = {2{`RANDOM}};
  tlb_sectored_entries_4_data_0 = _RAND_37[34:0];
  _RAND_38 = {2{`RANDOM}};
  tlb_sectored_entries_4_data_1 = _RAND_38[34:0];
  _RAND_39 = {2{`RANDOM}};
  tlb_sectored_entries_4_data_2 = _RAND_39[34:0];
  _RAND_40 = {2{`RANDOM}};
  tlb_sectored_entries_4_data_3 = _RAND_40[34:0];
  _RAND_41 = {1{`RANDOM}};
  tlb_sectored_entries_4_valid_0 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  tlb_sectored_entries_4_valid_1 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  tlb_sectored_entries_4_valid_2 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  tlb_sectored_entries_4_valid_3 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  tlb_sectored_entries_5_tag = _RAND_45[26:0];
  _RAND_46 = {2{`RANDOM}};
  tlb_sectored_entries_5_data_0 = _RAND_46[34:0];
  _RAND_47 = {2{`RANDOM}};
  tlb_sectored_entries_5_data_1 = _RAND_47[34:0];
  _RAND_48 = {2{`RANDOM}};
  tlb_sectored_entries_5_data_2 = _RAND_48[34:0];
  _RAND_49 = {2{`RANDOM}};
  tlb_sectored_entries_5_data_3 = _RAND_49[34:0];
  _RAND_50 = {1{`RANDOM}};
  tlb_sectored_entries_5_valid_0 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  tlb_sectored_entries_5_valid_1 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  tlb_sectored_entries_5_valid_2 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  tlb_sectored_entries_5_valid_3 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  tlb_sectored_entries_6_tag = _RAND_54[26:0];
  _RAND_55 = {2{`RANDOM}};
  tlb_sectored_entries_6_data_0 = _RAND_55[34:0];
  _RAND_56 = {2{`RANDOM}};
  tlb_sectored_entries_6_data_1 = _RAND_56[34:0];
  _RAND_57 = {2{`RANDOM}};
  tlb_sectored_entries_6_data_2 = _RAND_57[34:0];
  _RAND_58 = {2{`RANDOM}};
  tlb_sectored_entries_6_data_3 = _RAND_58[34:0];
  _RAND_59 = {1{`RANDOM}};
  tlb_sectored_entries_6_valid_0 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  tlb_sectored_entries_6_valid_1 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  tlb_sectored_entries_6_valid_2 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  tlb_sectored_entries_6_valid_3 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  tlb_sectored_entries_7_tag = _RAND_63[26:0];
  _RAND_64 = {2{`RANDOM}};
  tlb_sectored_entries_7_data_0 = _RAND_64[34:0];
  _RAND_65 = {2{`RANDOM}};
  tlb_sectored_entries_7_data_1 = _RAND_65[34:0];
  _RAND_66 = {2{`RANDOM}};
  tlb_sectored_entries_7_data_2 = _RAND_66[34:0];
  _RAND_67 = {2{`RANDOM}};
  tlb_sectored_entries_7_data_3 = _RAND_67[34:0];
  _RAND_68 = {1{`RANDOM}};
  tlb_sectored_entries_7_valid_0 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  tlb_sectored_entries_7_valid_1 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  tlb_sectored_entries_7_valid_2 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  tlb_sectored_entries_7_valid_3 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  tlb_superpage_entries_0_level = _RAND_72[1:0];
  _RAND_73 = {1{`RANDOM}};
  tlb_superpage_entries_0_tag = _RAND_73[26:0];
  _RAND_74 = {2{`RANDOM}};
  tlb_superpage_entries_0_data_0 = _RAND_74[34:0];
  _RAND_75 = {1{`RANDOM}};
  tlb_superpage_entries_0_valid_0 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  tlb_superpage_entries_1_level = _RAND_76[1:0];
  _RAND_77 = {1{`RANDOM}};
  tlb_superpage_entries_1_tag = _RAND_77[26:0];
  _RAND_78 = {2{`RANDOM}};
  tlb_superpage_entries_1_data_0 = _RAND_78[34:0];
  _RAND_79 = {1{`RANDOM}};
  tlb_superpage_entries_1_valid_0 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  tlb_superpage_entries_2_level = _RAND_80[1:0];
  _RAND_81 = {1{`RANDOM}};
  tlb_superpage_entries_2_tag = _RAND_81[26:0];
  _RAND_82 = {2{`RANDOM}};
  tlb_superpage_entries_2_data_0 = _RAND_82[34:0];
  _RAND_83 = {1{`RANDOM}};
  tlb_superpage_entries_2_valid_0 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  tlb_superpage_entries_3_level = _RAND_84[1:0];
  _RAND_85 = {1{`RANDOM}};
  tlb_superpage_entries_3_tag = _RAND_85[26:0];
  _RAND_86 = {2{`RANDOM}};
  tlb_superpage_entries_3_data_0 = _RAND_86[34:0];
  _RAND_87 = {1{`RANDOM}};
  tlb_superpage_entries_3_valid_0 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  tlb_special_entry_level = _RAND_88[1:0];
  _RAND_89 = {1{`RANDOM}};
  tlb_special_entry_tag = _RAND_89[26:0];
  _RAND_90 = {2{`RANDOM}};
  tlb_special_entry_data_0 = _RAND_90[34:0];
  _RAND_91 = {1{`RANDOM}};
  tlb_special_entry_valid_0 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  tlb_state = _RAND_92[1:0];
  _RAND_93 = {1{`RANDOM}};
  tlb_r_refill_tag = _RAND_93[26:0];
  _RAND_94 = {1{`RANDOM}};
  tlb_r_superpage_repl_addr = _RAND_94[1:0];
  _RAND_95 = {1{`RANDOM}};
  tlb_r_sectored_repl_addr = _RAND_95[2:0];
  _RAND_96 = {1{`RANDOM}};
  tlb_r_sectored_hit_addr = _RAND_96[2:0];
  _RAND_97 = {1{`RANDOM}};
  tlb_r_sectored_hit = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  tlb_state_reg = _RAND_98[6:0];
  _RAND_99 = {1{`RANDOM}};
  tlb_state_reg_1 = _RAND_99[2:0];
  _RAND_100 = {1{`RANDOM}};
  s1_valid = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  blockProbeAfterGrantCount = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  lrscCount = _RAND_102[6:0];
  _RAND_103 = {1{`RANDOM}};
  s1_probe = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  s2_probe = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  release_state = _RAND_105[2:0];
  _RAND_106 = {1{`RANDOM}};
  release_ack_wait = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  release_ack_addr = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  grantInProgress = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  s2_valid = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  probe_bits_param = _RAND_110[1:0];
  _RAND_111 = {1{`RANDOM}};
  probe_bits_size = _RAND_111[3:0];
  _RAND_112 = {1{`RANDOM}};
  probe_bits_source = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  probe_bits_address = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  s2_probe_state_state = _RAND_114[1:0];
  _RAND_115 = {1{`RANDOM}};
  counter_1 = _RAND_115[8:0];
  _RAND_116 = {1{`RANDOM}};
  s2_release_data_valid = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  s1_req_cmd = _RAND_117[4:0];
  _RAND_118 = {1{`RANDOM}};
  s2_req_cmd = _RAND_118[4:0];
  _RAND_119 = {1{`RANDOM}};
  pstore1_held = _RAND_119[0:0];
  _RAND_120 = {2{`RANDOM}};
  pstore1_addr = _RAND_120[39:0];
  _RAND_121 = {2{`RANDOM}};
  s1_req_addr = _RAND_121[39:0];
  _RAND_122 = {1{`RANDOM}};
  pstore1_mask = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  s1_req_size = _RAND_123[1:0];
  _RAND_124 = {1{`RANDOM}};
  pstore2_valid = _RAND_124[0:0];
  _RAND_125 = {2{`RANDOM}};
  pstore2_addr = _RAND_125[39:0];
  _RAND_126 = {1{`RANDOM}};
  mask = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  s2_not_nacked_in_s1 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  s2_hit_state_state = _RAND_128[1:0];
  _RAND_129 = {1{`RANDOM}};
  s1_req_tag = _RAND_129[6:0];
  _RAND_130 = {1{`RANDOM}};
  s1_req_signed = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  s1_req_dprv = _RAND_131[1:0];
  _RAND_132 = {2{`RANDOM}};
  s1_tlb_req_vaddr = _RAND_132[39:0];
  _RAND_133 = {1{`RANDOM}};
  s1_tlb_req_passthrough = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  s1_tlb_req_size = _RAND_134[1:0];
  _RAND_135 = {1{`RANDOM}};
  s1_tlb_req_cmd = _RAND_135[4:0];
  _RAND_136 = {1{`RANDOM}};
  cached_grant_wait = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  uncachedInFlight_0 = _RAND_137[0:0];
  _RAND_138 = {2{`RANDOM}};
  uncachedReqs_0_addr = _RAND_138[39:0];
  _RAND_139 = {1{`RANDOM}};
  uncachedReqs_0_tag = _RAND_139[6:0];
  _RAND_140 = {1{`RANDOM}};
  uncachedReqs_0_size = _RAND_140[1:0];
  _RAND_141 = {1{`RANDOM}};
  uncachedReqs_0_signed = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  s1_did_read = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  s2_hit_way = _RAND_143[3:0];
  _RAND_144 = {1{`RANDOM}};
  s2_victim_way_r = _RAND_144[1:0];
  _RAND_145 = {1{`RANDOM}};
  s2_probe_way = _RAND_145[3:0];
  _RAND_146 = {2{`RANDOM}};
  s2_req_addr = _RAND_146[39:0];
  _RAND_147 = {1{`RANDOM}};
  s2_req_tag = _RAND_147[6:0];
  _RAND_148 = {1{`RANDOM}};
  s2_req_size = _RAND_148[1:0];
  _RAND_149 = {1{`RANDOM}};
  s2_req_signed = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  s2_req_dprv = _RAND_150[1:0];
  _RAND_151 = {1{`RANDOM}};
  s2_tlb_xcpt_pf_ld = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  s2_tlb_xcpt_pf_st = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  s2_tlb_xcpt_ae_ld = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  s2_tlb_xcpt_ae_st = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  s2_tlb_xcpt_ma_ld = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  s2_tlb_xcpt_ma_st = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  s2_pma_cacheable = _RAND_157[0:0];
  _RAND_158 = {2{`RANDOM}};
  s2_uncached_resp_addr = _RAND_158[39:0];
  _RAND_159 = {2{`RANDOM}};
  s2_vaddr_r = _RAND_159[39:0];
  _RAND_160 = {1{`RANDOM}};
  blockUncachedGrant = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  counter = _RAND_161[8:0];
  _RAND_162 = {2{`RANDOM}};
  s2_data = _RAND_162[63:0];
  _RAND_163 = {1{`RANDOM}};
  s2_victim_tag_r = _RAND_163[19:0];
  _RAND_164 = {1{`RANDOM}};
  s2_victim_state_r_state = _RAND_164[1:0];
  _RAND_165 = {2{`RANDOM}};
  lrscAddr = _RAND_165[33:0];
  _RAND_166 = {1{`RANDOM}};
  pstore1_cmd = _RAND_166[4:0];
  _RAND_167 = {2{`RANDOM}};
  pstore1_data = _RAND_167[63:0];
  _RAND_168 = {1{`RANDOM}};
  pstore1_way = _RAND_168[3:0];
  _RAND_169 = {1{`RANDOM}};
  pstore1_rmw_r = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  pstore_drain_on_miss_REG = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  pstore2_way = _RAND_171[3:0];
  _RAND_172 = {1{`RANDOM}};
  pstore2_storegen_data_left_left_left = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  pstore2_storegen_data_left_left_right = _RAND_173[7:0];
  _RAND_174 = {1{`RANDOM}};
  pstore2_storegen_data_left_right_left = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  pstore2_storegen_data_left_right_right = _RAND_175[7:0];
  _RAND_176 = {1{`RANDOM}};
  pstore2_storegen_data_right_left_left = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  pstore2_storegen_data_right_left_right = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  pstore2_storegen_data_right_right_left = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  pstore2_storegen_data_right_right_right = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  s1_release_data_valid = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  io_cpu_s2_xcpt_REG = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  doUncachedResp = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  resetting = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  REG = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  flushCounter = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  io_cpu_perf_release_counter = _RAND_186[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
