module IntXbar(
  input   auto_int_in_0,
  input   auto_int_in_1,
  output  auto_int_out_0,
  output  auto_int_out_1
);
  assign auto_int_out_0 = auto_int_in_0; // @[Nodes.scala 1216:84 LazyModule.scala 312:16]
  assign auto_int_out_1 = auto_int_in_1; // @[Nodes.scala 1216:84 LazyModule.scala 312:16]
endmodule
