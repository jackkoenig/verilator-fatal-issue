module TLB_1(
  input         clock,
  input         reset,
  output        io_req_ready,
  input         io_req_valid,
  input  [39:0] io_req_bits_vaddr,
  output        io_resp_miss,
  output [31:0] io_resp_paddr,
  output        io_resp_pf_inst,
  output        io_resp_ae_inst,
  output        io_resp_cacheable,
  input         io_sfence_valid,
  input         io_sfence_bits_rs1,
  input         io_sfence_bits_rs2,
  input  [38:0] io_sfence_bits_addr,
  input         io_ptw_req_ready,
  output        io_ptw_req_valid,
  output        io_ptw_req_bits_valid,
  output [26:0] io_ptw_req_bits_bits_addr,
  input         io_ptw_resp_valid,
  input         io_ptw_resp_bits_ae,
  input  [53:0] io_ptw_resp_bits_pte_ppn,
  input         io_ptw_resp_bits_pte_d,
  input         io_ptw_resp_bits_pte_a,
  input         io_ptw_resp_bits_pte_g,
  input         io_ptw_resp_bits_pte_u,
  input         io_ptw_resp_bits_pte_x,
  input         io_ptw_resp_bits_pte_w,
  input         io_ptw_resp_bits_pte_r,
  input         io_ptw_resp_bits_pte_v,
  input  [1:0]  io_ptw_resp_bits_level,
  input         io_ptw_resp_bits_homogeneous,
  input  [3:0]  io_ptw_ptbr_mode,
  input         io_ptw_status_debug,
  input  [1:0]  io_ptw_status_prv,
  input         io_ptw_pmp_0_cfg_l,
  input  [1:0]  io_ptw_pmp_0_cfg_a,
  input         io_ptw_pmp_0_cfg_x,
  input         io_ptw_pmp_0_cfg_w,
  input         io_ptw_pmp_0_cfg_r,
  input  [29:0] io_ptw_pmp_0_addr,
  input  [31:0] io_ptw_pmp_0_mask,
  input         io_ptw_pmp_1_cfg_l,
  input  [1:0]  io_ptw_pmp_1_cfg_a,
  input         io_ptw_pmp_1_cfg_x,
  input         io_ptw_pmp_1_cfg_w,
  input         io_ptw_pmp_1_cfg_r,
  input  [29:0] io_ptw_pmp_1_addr,
  input  [31:0] io_ptw_pmp_1_mask,
  input         io_ptw_pmp_2_cfg_l,
  input  [1:0]  io_ptw_pmp_2_cfg_a,
  input         io_ptw_pmp_2_cfg_x,
  input         io_ptw_pmp_2_cfg_w,
  input         io_ptw_pmp_2_cfg_r,
  input  [29:0] io_ptw_pmp_2_addr,
  input  [31:0] io_ptw_pmp_2_mask,
  input         io_ptw_pmp_3_cfg_l,
  input  [1:0]  io_ptw_pmp_3_cfg_a,
  input         io_ptw_pmp_3_cfg_x,
  input         io_ptw_pmp_3_cfg_w,
  input         io_ptw_pmp_3_cfg_r,
  input  [29:0] io_ptw_pmp_3_addr,
  input  [31:0] io_ptw_pmp_3_mask,
  input         io_ptw_pmp_4_cfg_l,
  input  [1:0]  io_ptw_pmp_4_cfg_a,
  input         io_ptw_pmp_4_cfg_x,
  input         io_ptw_pmp_4_cfg_w,
  input         io_ptw_pmp_4_cfg_r,
  input  [29:0] io_ptw_pmp_4_addr,
  input  [31:0] io_ptw_pmp_4_mask,
  input         io_ptw_pmp_5_cfg_l,
  input  [1:0]  io_ptw_pmp_5_cfg_a,
  input         io_ptw_pmp_5_cfg_x,
  input         io_ptw_pmp_5_cfg_w,
  input         io_ptw_pmp_5_cfg_r,
  input  [29:0] io_ptw_pmp_5_addr,
  input  [31:0] io_ptw_pmp_5_mask,
  input         io_ptw_pmp_6_cfg_l,
  input  [1:0]  io_ptw_pmp_6_cfg_a,
  input         io_ptw_pmp_6_cfg_x,
  input         io_ptw_pmp_6_cfg_w,
  input         io_ptw_pmp_6_cfg_r,
  input  [29:0] io_ptw_pmp_6_addr,
  input  [31:0] io_ptw_pmp_6_mask,
  input         io_ptw_pmp_7_cfg_l,
  input  [1:0]  io_ptw_pmp_7_cfg_a,
  input         io_ptw_pmp_7_cfg_x,
  input         io_ptw_pmp_7_cfg_w,
  input         io_ptw_pmp_7_cfg_r,
  input  [29:0] io_ptw_pmp_7_addr,
  input  [31:0] io_ptw_pmp_7_mask,
  input         io_kill
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [63:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
`endif // RANDOMIZE_REG_INIT
  wire [19:0] mpu_ppn_data_barrier_io_x_ppn; // @[package.scala 236:25]
  wire  mpu_ppn_data_barrier_io_x_u; // @[package.scala 236:25]
  wire  mpu_ppn_data_barrier_io_x_ae; // @[package.scala 236:25]
  wire  mpu_ppn_data_barrier_io_x_sw; // @[package.scala 236:25]
  wire  mpu_ppn_data_barrier_io_x_sx; // @[package.scala 236:25]
  wire  mpu_ppn_data_barrier_io_x_sr; // @[package.scala 236:25]
  wire  mpu_ppn_data_barrier_io_x_pw; // @[package.scala 236:25]
  wire  mpu_ppn_data_barrier_io_x_px; // @[package.scala 236:25]
  wire  mpu_ppn_data_barrier_io_x_pr; // @[package.scala 236:25]
  wire  mpu_ppn_data_barrier_io_x_ppp; // @[package.scala 236:25]
  wire  mpu_ppn_data_barrier_io_x_pal; // @[package.scala 236:25]
  wire  mpu_ppn_data_barrier_io_x_paa; // @[package.scala 236:25]
  wire  mpu_ppn_data_barrier_io_x_eff; // @[package.scala 236:25]
  wire  mpu_ppn_data_barrier_io_x_c; // @[package.scala 236:25]
  wire [19:0] mpu_ppn_data_barrier_io_y_ppn; // @[package.scala 236:25]
  wire  mpu_ppn_data_barrier_io_y_u; // @[package.scala 236:25]
  wire  mpu_ppn_data_barrier_io_y_ae; // @[package.scala 236:25]
  wire  mpu_ppn_data_barrier_io_y_sw; // @[package.scala 236:25]
  wire  mpu_ppn_data_barrier_io_y_sx; // @[package.scala 236:25]
  wire  mpu_ppn_data_barrier_io_y_sr; // @[package.scala 236:25]
  wire  mpu_ppn_data_barrier_io_y_pw; // @[package.scala 236:25]
  wire  mpu_ppn_data_barrier_io_y_px; // @[package.scala 236:25]
  wire  mpu_ppn_data_barrier_io_y_pr; // @[package.scala 236:25]
  wire  mpu_ppn_data_barrier_io_y_ppp; // @[package.scala 236:25]
  wire  mpu_ppn_data_barrier_io_y_pal; // @[package.scala 236:25]
  wire  mpu_ppn_data_barrier_io_y_paa; // @[package.scala 236:25]
  wire  mpu_ppn_data_barrier_io_y_eff; // @[package.scala 236:25]
  wire  mpu_ppn_data_barrier_io_y_c; // @[package.scala 236:25]
  wire [1:0] pmp_io_prv; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_0_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_0_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_0_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_0_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_0_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_0_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_0_mask; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_1_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_1_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_1_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_1_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_1_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_1_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_1_mask; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_2_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_2_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_2_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_2_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_2_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_2_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_2_mask; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_3_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_3_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_3_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_3_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_3_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_3_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_3_mask; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_4_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_4_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_4_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_4_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_4_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_4_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_4_mask; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_5_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_5_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_5_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_5_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_5_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_5_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_5_mask; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_6_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_6_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_6_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_6_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_6_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_6_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_6_mask; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_7_cfg_l; // @[TLB.scala 190:19]
  wire [1:0] pmp_io_pmp_7_cfg_a; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_7_cfg_x; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_7_cfg_w; // @[TLB.scala 190:19]
  wire  pmp_io_pmp_7_cfg_r; // @[TLB.scala 190:19]
  wire [29:0] pmp_io_pmp_7_addr; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_pmp_7_mask; // @[TLB.scala 190:19]
  wire [31:0] pmp_io_addr; // @[TLB.scala 190:19]
  wire  pmp_io_r; // @[TLB.scala 190:19]
  wire  pmp_io_w; // @[TLB.scala 190:19]
  wire  pmp_io_x; // @[TLB.scala 190:19]
  wire [19:0] ppn_data_barrier_io_x_ppn; // @[package.scala 236:25]
  wire  ppn_data_barrier_io_x_u; // @[package.scala 236:25]
  wire  ppn_data_barrier_io_x_ae; // @[package.scala 236:25]
  wire  ppn_data_barrier_io_x_sw; // @[package.scala 236:25]
  wire  ppn_data_barrier_io_x_sx; // @[package.scala 236:25]
  wire  ppn_data_barrier_io_x_sr; // @[package.scala 236:25]
  wire  ppn_data_barrier_io_x_pw; // @[package.scala 236:25]
  wire  ppn_data_barrier_io_x_px; // @[package.scala 236:25]
  wire  ppn_data_barrier_io_x_pr; // @[package.scala 236:25]
  wire  ppn_data_barrier_io_x_ppp; // @[package.scala 236:25]
  wire  ppn_data_barrier_io_x_pal; // @[package.scala 236:25]
  wire  ppn_data_barrier_io_x_paa; // @[package.scala 236:25]
  wire  ppn_data_barrier_io_x_eff; // @[package.scala 236:25]
  wire  ppn_data_barrier_io_x_c; // @[package.scala 236:25]
  wire [19:0] ppn_data_barrier_io_y_ppn; // @[package.scala 236:25]
  wire  ppn_data_barrier_io_y_u; // @[package.scala 236:25]
  wire  ppn_data_barrier_io_y_ae; // @[package.scala 236:25]
  wire  ppn_data_barrier_io_y_sw; // @[package.scala 236:25]
  wire  ppn_data_barrier_io_y_sx; // @[package.scala 236:25]
  wire  ppn_data_barrier_io_y_sr; // @[package.scala 236:25]
  wire  ppn_data_barrier_io_y_pw; // @[package.scala 236:25]
  wire  ppn_data_barrier_io_y_px; // @[package.scala 236:25]
  wire  ppn_data_barrier_io_y_pr; // @[package.scala 236:25]
  wire  ppn_data_barrier_io_y_ppp; // @[package.scala 236:25]
  wire  ppn_data_barrier_io_y_pal; // @[package.scala 236:25]
  wire  ppn_data_barrier_io_y_paa; // @[package.scala 236:25]
  wire  ppn_data_barrier_io_y_eff; // @[package.scala 236:25]
  wire  ppn_data_barrier_io_y_c; // @[package.scala 236:25]
  wire [19:0] ppn_data_barrier_1_io_x_ppn; // @[package.scala 236:25]
  wire  ppn_data_barrier_1_io_x_u; // @[package.scala 236:25]
  wire  ppn_data_barrier_1_io_x_ae; // @[package.scala 236:25]
  wire  ppn_data_barrier_1_io_x_sw; // @[package.scala 236:25]
  wire  ppn_data_barrier_1_io_x_sx; // @[package.scala 236:25]
  wire  ppn_data_barrier_1_io_x_sr; // @[package.scala 236:25]
  wire  ppn_data_barrier_1_io_x_pw; // @[package.scala 236:25]
  wire  ppn_data_barrier_1_io_x_px; // @[package.scala 236:25]
  wire  ppn_data_barrier_1_io_x_pr; // @[package.scala 236:25]
  wire  ppn_data_barrier_1_io_x_ppp; // @[package.scala 236:25]
  wire  ppn_data_barrier_1_io_x_pal; // @[package.scala 236:25]
  wire  ppn_data_barrier_1_io_x_paa; // @[package.scala 236:25]
  wire  ppn_data_barrier_1_io_x_eff; // @[package.scala 236:25]
  wire  ppn_data_barrier_1_io_x_c; // @[package.scala 236:25]
  wire [19:0] ppn_data_barrier_1_io_y_ppn; // @[package.scala 236:25]
  wire  ppn_data_barrier_1_io_y_u; // @[package.scala 236:25]
  wire  ppn_data_barrier_1_io_y_ae; // @[package.scala 236:25]
  wire  ppn_data_barrier_1_io_y_sw; // @[package.scala 236:25]
  wire  ppn_data_barrier_1_io_y_sx; // @[package.scala 236:25]
  wire  ppn_data_barrier_1_io_y_sr; // @[package.scala 236:25]
  wire  ppn_data_barrier_1_io_y_pw; // @[package.scala 236:25]
  wire  ppn_data_barrier_1_io_y_px; // @[package.scala 236:25]
  wire  ppn_data_barrier_1_io_y_pr; // @[package.scala 236:25]
  wire  ppn_data_barrier_1_io_y_ppp; // @[package.scala 236:25]
  wire  ppn_data_barrier_1_io_y_pal; // @[package.scala 236:25]
  wire  ppn_data_barrier_1_io_y_paa; // @[package.scala 236:25]
  wire  ppn_data_barrier_1_io_y_eff; // @[package.scala 236:25]
  wire  ppn_data_barrier_1_io_y_c; // @[package.scala 236:25]
  wire [19:0] ppn_data_barrier_2_io_x_ppn; // @[package.scala 236:25]
  wire  ppn_data_barrier_2_io_x_u; // @[package.scala 236:25]
  wire  ppn_data_barrier_2_io_x_ae; // @[package.scala 236:25]
  wire  ppn_data_barrier_2_io_x_sw; // @[package.scala 236:25]
  wire  ppn_data_barrier_2_io_x_sx; // @[package.scala 236:25]
  wire  ppn_data_barrier_2_io_x_sr; // @[package.scala 236:25]
  wire  ppn_data_barrier_2_io_x_pw; // @[package.scala 236:25]
  wire  ppn_data_barrier_2_io_x_px; // @[package.scala 236:25]
  wire  ppn_data_barrier_2_io_x_pr; // @[package.scala 236:25]
  wire  ppn_data_barrier_2_io_x_ppp; // @[package.scala 236:25]
  wire  ppn_data_barrier_2_io_x_pal; // @[package.scala 236:25]
  wire  ppn_data_barrier_2_io_x_paa; // @[package.scala 236:25]
  wire  ppn_data_barrier_2_io_x_eff; // @[package.scala 236:25]
  wire  ppn_data_barrier_2_io_x_c; // @[package.scala 236:25]
  wire [19:0] ppn_data_barrier_2_io_y_ppn; // @[package.scala 236:25]
  wire  ppn_data_barrier_2_io_y_u; // @[package.scala 236:25]
  wire  ppn_data_barrier_2_io_y_ae; // @[package.scala 236:25]
  wire  ppn_data_barrier_2_io_y_sw; // @[package.scala 236:25]
  wire  ppn_data_barrier_2_io_y_sx; // @[package.scala 236:25]
  wire  ppn_data_barrier_2_io_y_sr; // @[package.scala 236:25]
  wire  ppn_data_barrier_2_io_y_pw; // @[package.scala 236:25]
  wire  ppn_data_barrier_2_io_y_px; // @[package.scala 236:25]
  wire  ppn_data_barrier_2_io_y_pr; // @[package.scala 236:25]
  wire  ppn_data_barrier_2_io_y_ppp; // @[package.scala 236:25]
  wire  ppn_data_barrier_2_io_y_pal; // @[package.scala 236:25]
  wire  ppn_data_barrier_2_io_y_paa; // @[package.scala 236:25]
  wire  ppn_data_barrier_2_io_y_eff; // @[package.scala 236:25]
  wire  ppn_data_barrier_2_io_y_c; // @[package.scala 236:25]
  wire [19:0] ppn_data_barrier_3_io_x_ppn; // @[package.scala 236:25]
  wire  ppn_data_barrier_3_io_x_u; // @[package.scala 236:25]
  wire  ppn_data_barrier_3_io_x_ae; // @[package.scala 236:25]
  wire  ppn_data_barrier_3_io_x_sw; // @[package.scala 236:25]
  wire  ppn_data_barrier_3_io_x_sx; // @[package.scala 236:25]
  wire  ppn_data_barrier_3_io_x_sr; // @[package.scala 236:25]
  wire  ppn_data_barrier_3_io_x_pw; // @[package.scala 236:25]
  wire  ppn_data_barrier_3_io_x_px; // @[package.scala 236:25]
  wire  ppn_data_barrier_3_io_x_pr; // @[package.scala 236:25]
  wire  ppn_data_barrier_3_io_x_ppp; // @[package.scala 236:25]
  wire  ppn_data_barrier_3_io_x_pal; // @[package.scala 236:25]
  wire  ppn_data_barrier_3_io_x_paa; // @[package.scala 236:25]
  wire  ppn_data_barrier_3_io_x_eff; // @[package.scala 236:25]
  wire  ppn_data_barrier_3_io_x_c; // @[package.scala 236:25]
  wire [19:0] ppn_data_barrier_3_io_y_ppn; // @[package.scala 236:25]
  wire  ppn_data_barrier_3_io_y_u; // @[package.scala 236:25]
  wire  ppn_data_barrier_3_io_y_ae; // @[package.scala 236:25]
  wire  ppn_data_barrier_3_io_y_sw; // @[package.scala 236:25]
  wire  ppn_data_barrier_3_io_y_sx; // @[package.scala 236:25]
  wire  ppn_data_barrier_3_io_y_sr; // @[package.scala 236:25]
  wire  ppn_data_barrier_3_io_y_pw; // @[package.scala 236:25]
  wire  ppn_data_barrier_3_io_y_px; // @[package.scala 236:25]
  wire  ppn_data_barrier_3_io_y_pr; // @[package.scala 236:25]
  wire  ppn_data_barrier_3_io_y_ppp; // @[package.scala 236:25]
  wire  ppn_data_barrier_3_io_y_pal; // @[package.scala 236:25]
  wire  ppn_data_barrier_3_io_y_paa; // @[package.scala 236:25]
  wire  ppn_data_barrier_3_io_y_eff; // @[package.scala 236:25]
  wire  ppn_data_barrier_3_io_y_c; // @[package.scala 236:25]
  wire [19:0] ppn_data_barrier_4_io_x_ppn; // @[package.scala 236:25]
  wire  ppn_data_barrier_4_io_x_u; // @[package.scala 236:25]
  wire  ppn_data_barrier_4_io_x_ae; // @[package.scala 236:25]
  wire  ppn_data_barrier_4_io_x_sw; // @[package.scala 236:25]
  wire  ppn_data_barrier_4_io_x_sx; // @[package.scala 236:25]
  wire  ppn_data_barrier_4_io_x_sr; // @[package.scala 236:25]
  wire  ppn_data_barrier_4_io_x_pw; // @[package.scala 236:25]
  wire  ppn_data_barrier_4_io_x_px; // @[package.scala 236:25]
  wire  ppn_data_barrier_4_io_x_pr; // @[package.scala 236:25]
  wire  ppn_data_barrier_4_io_x_ppp; // @[package.scala 236:25]
  wire  ppn_data_barrier_4_io_x_pal; // @[package.scala 236:25]
  wire  ppn_data_barrier_4_io_x_paa; // @[package.scala 236:25]
  wire  ppn_data_barrier_4_io_x_eff; // @[package.scala 236:25]
  wire  ppn_data_barrier_4_io_x_c; // @[package.scala 236:25]
  wire [19:0] ppn_data_barrier_4_io_y_ppn; // @[package.scala 236:25]
  wire  ppn_data_barrier_4_io_y_u; // @[package.scala 236:25]
  wire  ppn_data_barrier_4_io_y_ae; // @[package.scala 236:25]
  wire  ppn_data_barrier_4_io_y_sw; // @[package.scala 236:25]
  wire  ppn_data_barrier_4_io_y_sx; // @[package.scala 236:25]
  wire  ppn_data_barrier_4_io_y_sr; // @[package.scala 236:25]
  wire  ppn_data_barrier_4_io_y_pw; // @[package.scala 236:25]
  wire  ppn_data_barrier_4_io_y_px; // @[package.scala 236:25]
  wire  ppn_data_barrier_4_io_y_pr; // @[package.scala 236:25]
  wire  ppn_data_barrier_4_io_y_ppp; // @[package.scala 236:25]
  wire  ppn_data_barrier_4_io_y_pal; // @[package.scala 236:25]
  wire  ppn_data_barrier_4_io_y_paa; // @[package.scala 236:25]
  wire  ppn_data_barrier_4_io_y_eff; // @[package.scala 236:25]
  wire  ppn_data_barrier_4_io_y_c; // @[package.scala 236:25]
  wire [19:0] ppn_data_barrier_5_io_x_ppn; // @[package.scala 236:25]
  wire  ppn_data_barrier_5_io_x_u; // @[package.scala 236:25]
  wire  ppn_data_barrier_5_io_x_ae; // @[package.scala 236:25]
  wire  ppn_data_barrier_5_io_x_sw; // @[package.scala 236:25]
  wire  ppn_data_barrier_5_io_x_sx; // @[package.scala 236:25]
  wire  ppn_data_barrier_5_io_x_sr; // @[package.scala 236:25]
  wire  ppn_data_barrier_5_io_x_pw; // @[package.scala 236:25]
  wire  ppn_data_barrier_5_io_x_px; // @[package.scala 236:25]
  wire  ppn_data_barrier_5_io_x_pr; // @[package.scala 236:25]
  wire  ppn_data_barrier_5_io_x_ppp; // @[package.scala 236:25]
  wire  ppn_data_barrier_5_io_x_pal; // @[package.scala 236:25]
  wire  ppn_data_barrier_5_io_x_paa; // @[package.scala 236:25]
  wire  ppn_data_barrier_5_io_x_eff; // @[package.scala 236:25]
  wire  ppn_data_barrier_5_io_x_c; // @[package.scala 236:25]
  wire [19:0] ppn_data_barrier_5_io_y_ppn; // @[package.scala 236:25]
  wire  ppn_data_barrier_5_io_y_u; // @[package.scala 236:25]
  wire  ppn_data_barrier_5_io_y_ae; // @[package.scala 236:25]
  wire  ppn_data_barrier_5_io_y_sw; // @[package.scala 236:25]
  wire  ppn_data_barrier_5_io_y_sx; // @[package.scala 236:25]
  wire  ppn_data_barrier_5_io_y_sr; // @[package.scala 236:25]
  wire  ppn_data_barrier_5_io_y_pw; // @[package.scala 236:25]
  wire  ppn_data_barrier_5_io_y_px; // @[package.scala 236:25]
  wire  ppn_data_barrier_5_io_y_pr; // @[package.scala 236:25]
  wire  ppn_data_barrier_5_io_y_ppp; // @[package.scala 236:25]
  wire  ppn_data_barrier_5_io_y_pal; // @[package.scala 236:25]
  wire  ppn_data_barrier_5_io_y_paa; // @[package.scala 236:25]
  wire  ppn_data_barrier_5_io_y_eff; // @[package.scala 236:25]
  wire  ppn_data_barrier_5_io_y_c; // @[package.scala 236:25]
  wire [19:0] ppn_data_barrier_6_io_x_ppn; // @[package.scala 236:25]
  wire  ppn_data_barrier_6_io_x_u; // @[package.scala 236:25]
  wire  ppn_data_barrier_6_io_x_ae; // @[package.scala 236:25]
  wire  ppn_data_barrier_6_io_x_sw; // @[package.scala 236:25]
  wire  ppn_data_barrier_6_io_x_sx; // @[package.scala 236:25]
  wire  ppn_data_barrier_6_io_x_sr; // @[package.scala 236:25]
  wire  ppn_data_barrier_6_io_x_pw; // @[package.scala 236:25]
  wire  ppn_data_barrier_6_io_x_px; // @[package.scala 236:25]
  wire  ppn_data_barrier_6_io_x_pr; // @[package.scala 236:25]
  wire  ppn_data_barrier_6_io_x_ppp; // @[package.scala 236:25]
  wire  ppn_data_barrier_6_io_x_pal; // @[package.scala 236:25]
  wire  ppn_data_barrier_6_io_x_paa; // @[package.scala 236:25]
  wire  ppn_data_barrier_6_io_x_eff; // @[package.scala 236:25]
  wire  ppn_data_barrier_6_io_x_c; // @[package.scala 236:25]
  wire [19:0] ppn_data_barrier_6_io_y_ppn; // @[package.scala 236:25]
  wire  ppn_data_barrier_6_io_y_u; // @[package.scala 236:25]
  wire  ppn_data_barrier_6_io_y_ae; // @[package.scala 236:25]
  wire  ppn_data_barrier_6_io_y_sw; // @[package.scala 236:25]
  wire  ppn_data_barrier_6_io_y_sx; // @[package.scala 236:25]
  wire  ppn_data_barrier_6_io_y_sr; // @[package.scala 236:25]
  wire  ppn_data_barrier_6_io_y_pw; // @[package.scala 236:25]
  wire  ppn_data_barrier_6_io_y_px; // @[package.scala 236:25]
  wire  ppn_data_barrier_6_io_y_pr; // @[package.scala 236:25]
  wire  ppn_data_barrier_6_io_y_ppp; // @[package.scala 236:25]
  wire  ppn_data_barrier_6_io_y_pal; // @[package.scala 236:25]
  wire  ppn_data_barrier_6_io_y_paa; // @[package.scala 236:25]
  wire  ppn_data_barrier_6_io_y_eff; // @[package.scala 236:25]
  wire  ppn_data_barrier_6_io_y_c; // @[package.scala 236:25]
  wire [19:0] ppn_data_barrier_7_io_x_ppn; // @[package.scala 236:25]
  wire  ppn_data_barrier_7_io_x_u; // @[package.scala 236:25]
  wire  ppn_data_barrier_7_io_x_ae; // @[package.scala 236:25]
  wire  ppn_data_barrier_7_io_x_sw; // @[package.scala 236:25]
  wire  ppn_data_barrier_7_io_x_sx; // @[package.scala 236:25]
  wire  ppn_data_barrier_7_io_x_sr; // @[package.scala 236:25]
  wire  ppn_data_barrier_7_io_x_pw; // @[package.scala 236:25]
  wire  ppn_data_barrier_7_io_x_px; // @[package.scala 236:25]
  wire  ppn_data_barrier_7_io_x_pr; // @[package.scala 236:25]
  wire  ppn_data_barrier_7_io_x_ppp; // @[package.scala 236:25]
  wire  ppn_data_barrier_7_io_x_pal; // @[package.scala 236:25]
  wire  ppn_data_barrier_7_io_x_paa; // @[package.scala 236:25]
  wire  ppn_data_barrier_7_io_x_eff; // @[package.scala 236:25]
  wire  ppn_data_barrier_7_io_x_c; // @[package.scala 236:25]
  wire [19:0] ppn_data_barrier_7_io_y_ppn; // @[package.scala 236:25]
  wire  ppn_data_barrier_7_io_y_u; // @[package.scala 236:25]
  wire  ppn_data_barrier_7_io_y_ae; // @[package.scala 236:25]
  wire  ppn_data_barrier_7_io_y_sw; // @[package.scala 236:25]
  wire  ppn_data_barrier_7_io_y_sx; // @[package.scala 236:25]
  wire  ppn_data_barrier_7_io_y_sr; // @[package.scala 236:25]
  wire  ppn_data_barrier_7_io_y_pw; // @[package.scala 236:25]
  wire  ppn_data_barrier_7_io_y_px; // @[package.scala 236:25]
  wire  ppn_data_barrier_7_io_y_pr; // @[package.scala 236:25]
  wire  ppn_data_barrier_7_io_y_ppp; // @[package.scala 236:25]
  wire  ppn_data_barrier_7_io_y_pal; // @[package.scala 236:25]
  wire  ppn_data_barrier_7_io_y_paa; // @[package.scala 236:25]
  wire  ppn_data_barrier_7_io_y_eff; // @[package.scala 236:25]
  wire  ppn_data_barrier_7_io_y_c; // @[package.scala 236:25]
  wire [19:0] ppn_data_barrier_8_io_x_ppn; // @[package.scala 236:25]
  wire  ppn_data_barrier_8_io_x_u; // @[package.scala 236:25]
  wire  ppn_data_barrier_8_io_x_ae; // @[package.scala 236:25]
  wire  ppn_data_barrier_8_io_x_sw; // @[package.scala 236:25]
  wire  ppn_data_barrier_8_io_x_sx; // @[package.scala 236:25]
  wire  ppn_data_barrier_8_io_x_sr; // @[package.scala 236:25]
  wire  ppn_data_barrier_8_io_x_pw; // @[package.scala 236:25]
  wire  ppn_data_barrier_8_io_x_px; // @[package.scala 236:25]
  wire  ppn_data_barrier_8_io_x_pr; // @[package.scala 236:25]
  wire  ppn_data_barrier_8_io_x_ppp; // @[package.scala 236:25]
  wire  ppn_data_barrier_8_io_x_pal; // @[package.scala 236:25]
  wire  ppn_data_barrier_8_io_x_paa; // @[package.scala 236:25]
  wire  ppn_data_barrier_8_io_x_eff; // @[package.scala 236:25]
  wire  ppn_data_barrier_8_io_x_c; // @[package.scala 236:25]
  wire [19:0] ppn_data_barrier_8_io_y_ppn; // @[package.scala 236:25]
  wire  ppn_data_barrier_8_io_y_u; // @[package.scala 236:25]
  wire  ppn_data_barrier_8_io_y_ae; // @[package.scala 236:25]
  wire  ppn_data_barrier_8_io_y_sw; // @[package.scala 236:25]
  wire  ppn_data_barrier_8_io_y_sx; // @[package.scala 236:25]
  wire  ppn_data_barrier_8_io_y_sr; // @[package.scala 236:25]
  wire  ppn_data_barrier_8_io_y_pw; // @[package.scala 236:25]
  wire  ppn_data_barrier_8_io_y_px; // @[package.scala 236:25]
  wire  ppn_data_barrier_8_io_y_pr; // @[package.scala 236:25]
  wire  ppn_data_barrier_8_io_y_ppp; // @[package.scala 236:25]
  wire  ppn_data_barrier_8_io_y_pal; // @[package.scala 236:25]
  wire  ppn_data_barrier_8_io_y_paa; // @[package.scala 236:25]
  wire  ppn_data_barrier_8_io_y_eff; // @[package.scala 236:25]
  wire  ppn_data_barrier_8_io_y_c; // @[package.scala 236:25]
  wire [19:0] ppn_data_barrier_9_io_x_ppn; // @[package.scala 236:25]
  wire  ppn_data_barrier_9_io_x_u; // @[package.scala 236:25]
  wire  ppn_data_barrier_9_io_x_ae; // @[package.scala 236:25]
  wire  ppn_data_barrier_9_io_x_sw; // @[package.scala 236:25]
  wire  ppn_data_barrier_9_io_x_sx; // @[package.scala 236:25]
  wire  ppn_data_barrier_9_io_x_sr; // @[package.scala 236:25]
  wire  ppn_data_barrier_9_io_x_pw; // @[package.scala 236:25]
  wire  ppn_data_barrier_9_io_x_px; // @[package.scala 236:25]
  wire  ppn_data_barrier_9_io_x_pr; // @[package.scala 236:25]
  wire  ppn_data_barrier_9_io_x_ppp; // @[package.scala 236:25]
  wire  ppn_data_barrier_9_io_x_pal; // @[package.scala 236:25]
  wire  ppn_data_barrier_9_io_x_paa; // @[package.scala 236:25]
  wire  ppn_data_barrier_9_io_x_eff; // @[package.scala 236:25]
  wire  ppn_data_barrier_9_io_x_c; // @[package.scala 236:25]
  wire [19:0] ppn_data_barrier_9_io_y_ppn; // @[package.scala 236:25]
  wire  ppn_data_barrier_9_io_y_u; // @[package.scala 236:25]
  wire  ppn_data_barrier_9_io_y_ae; // @[package.scala 236:25]
  wire  ppn_data_barrier_9_io_y_sw; // @[package.scala 236:25]
  wire  ppn_data_barrier_9_io_y_sx; // @[package.scala 236:25]
  wire  ppn_data_barrier_9_io_y_sr; // @[package.scala 236:25]
  wire  ppn_data_barrier_9_io_y_pw; // @[package.scala 236:25]
  wire  ppn_data_barrier_9_io_y_px; // @[package.scala 236:25]
  wire  ppn_data_barrier_9_io_y_pr; // @[package.scala 236:25]
  wire  ppn_data_barrier_9_io_y_ppp; // @[package.scala 236:25]
  wire  ppn_data_barrier_9_io_y_pal; // @[package.scala 236:25]
  wire  ppn_data_barrier_9_io_y_paa; // @[package.scala 236:25]
  wire  ppn_data_barrier_9_io_y_eff; // @[package.scala 236:25]
  wire  ppn_data_barrier_9_io_y_c; // @[package.scala 236:25]
  wire [19:0] ppn_data_barrier_10_io_x_ppn; // @[package.scala 236:25]
  wire  ppn_data_barrier_10_io_x_u; // @[package.scala 236:25]
  wire  ppn_data_barrier_10_io_x_ae; // @[package.scala 236:25]
  wire  ppn_data_barrier_10_io_x_sw; // @[package.scala 236:25]
  wire  ppn_data_barrier_10_io_x_sx; // @[package.scala 236:25]
  wire  ppn_data_barrier_10_io_x_sr; // @[package.scala 236:25]
  wire  ppn_data_barrier_10_io_x_pw; // @[package.scala 236:25]
  wire  ppn_data_barrier_10_io_x_px; // @[package.scala 236:25]
  wire  ppn_data_barrier_10_io_x_pr; // @[package.scala 236:25]
  wire  ppn_data_barrier_10_io_x_ppp; // @[package.scala 236:25]
  wire  ppn_data_barrier_10_io_x_pal; // @[package.scala 236:25]
  wire  ppn_data_barrier_10_io_x_paa; // @[package.scala 236:25]
  wire  ppn_data_barrier_10_io_x_eff; // @[package.scala 236:25]
  wire  ppn_data_barrier_10_io_x_c; // @[package.scala 236:25]
  wire [19:0] ppn_data_barrier_10_io_y_ppn; // @[package.scala 236:25]
  wire  ppn_data_barrier_10_io_y_u; // @[package.scala 236:25]
  wire  ppn_data_barrier_10_io_y_ae; // @[package.scala 236:25]
  wire  ppn_data_barrier_10_io_y_sw; // @[package.scala 236:25]
  wire  ppn_data_barrier_10_io_y_sx; // @[package.scala 236:25]
  wire  ppn_data_barrier_10_io_y_sr; // @[package.scala 236:25]
  wire  ppn_data_barrier_10_io_y_pw; // @[package.scala 236:25]
  wire  ppn_data_barrier_10_io_y_px; // @[package.scala 236:25]
  wire  ppn_data_barrier_10_io_y_pr; // @[package.scala 236:25]
  wire  ppn_data_barrier_10_io_y_ppp; // @[package.scala 236:25]
  wire  ppn_data_barrier_10_io_y_pal; // @[package.scala 236:25]
  wire  ppn_data_barrier_10_io_y_paa; // @[package.scala 236:25]
  wire  ppn_data_barrier_10_io_y_eff; // @[package.scala 236:25]
  wire  ppn_data_barrier_10_io_y_c; // @[package.scala 236:25]
  wire [19:0] ppn_data_barrier_11_io_x_ppn; // @[package.scala 236:25]
  wire  ppn_data_barrier_11_io_x_u; // @[package.scala 236:25]
  wire  ppn_data_barrier_11_io_x_ae; // @[package.scala 236:25]
  wire  ppn_data_barrier_11_io_x_sw; // @[package.scala 236:25]
  wire  ppn_data_barrier_11_io_x_sx; // @[package.scala 236:25]
  wire  ppn_data_barrier_11_io_x_sr; // @[package.scala 236:25]
  wire  ppn_data_barrier_11_io_x_pw; // @[package.scala 236:25]
  wire  ppn_data_barrier_11_io_x_px; // @[package.scala 236:25]
  wire  ppn_data_barrier_11_io_x_pr; // @[package.scala 236:25]
  wire  ppn_data_barrier_11_io_x_ppp; // @[package.scala 236:25]
  wire  ppn_data_barrier_11_io_x_pal; // @[package.scala 236:25]
  wire  ppn_data_barrier_11_io_x_paa; // @[package.scala 236:25]
  wire  ppn_data_barrier_11_io_x_eff; // @[package.scala 236:25]
  wire  ppn_data_barrier_11_io_x_c; // @[package.scala 236:25]
  wire [19:0] ppn_data_barrier_11_io_y_ppn; // @[package.scala 236:25]
  wire  ppn_data_barrier_11_io_y_u; // @[package.scala 236:25]
  wire  ppn_data_barrier_11_io_y_ae; // @[package.scala 236:25]
  wire  ppn_data_barrier_11_io_y_sw; // @[package.scala 236:25]
  wire  ppn_data_barrier_11_io_y_sx; // @[package.scala 236:25]
  wire  ppn_data_barrier_11_io_y_sr; // @[package.scala 236:25]
  wire  ppn_data_barrier_11_io_y_pw; // @[package.scala 236:25]
  wire  ppn_data_barrier_11_io_y_px; // @[package.scala 236:25]
  wire  ppn_data_barrier_11_io_y_pr; // @[package.scala 236:25]
  wire  ppn_data_barrier_11_io_y_ppp; // @[package.scala 236:25]
  wire  ppn_data_barrier_11_io_y_pal; // @[package.scala 236:25]
  wire  ppn_data_barrier_11_io_y_paa; // @[package.scala 236:25]
  wire  ppn_data_barrier_11_io_y_eff; // @[package.scala 236:25]
  wire  ppn_data_barrier_11_io_y_c; // @[package.scala 236:25]
  wire [19:0] ppn_data_barrier_12_io_x_ppn; // @[package.scala 236:25]
  wire  ppn_data_barrier_12_io_x_u; // @[package.scala 236:25]
  wire  ppn_data_barrier_12_io_x_ae; // @[package.scala 236:25]
  wire  ppn_data_barrier_12_io_x_sw; // @[package.scala 236:25]
  wire  ppn_data_barrier_12_io_x_sx; // @[package.scala 236:25]
  wire  ppn_data_barrier_12_io_x_sr; // @[package.scala 236:25]
  wire  ppn_data_barrier_12_io_x_pw; // @[package.scala 236:25]
  wire  ppn_data_barrier_12_io_x_px; // @[package.scala 236:25]
  wire  ppn_data_barrier_12_io_x_pr; // @[package.scala 236:25]
  wire  ppn_data_barrier_12_io_x_ppp; // @[package.scala 236:25]
  wire  ppn_data_barrier_12_io_x_pal; // @[package.scala 236:25]
  wire  ppn_data_barrier_12_io_x_paa; // @[package.scala 236:25]
  wire  ppn_data_barrier_12_io_x_eff; // @[package.scala 236:25]
  wire  ppn_data_barrier_12_io_x_c; // @[package.scala 236:25]
  wire [19:0] ppn_data_barrier_12_io_y_ppn; // @[package.scala 236:25]
  wire  ppn_data_barrier_12_io_y_u; // @[package.scala 236:25]
  wire  ppn_data_barrier_12_io_y_ae; // @[package.scala 236:25]
  wire  ppn_data_barrier_12_io_y_sw; // @[package.scala 236:25]
  wire  ppn_data_barrier_12_io_y_sx; // @[package.scala 236:25]
  wire  ppn_data_barrier_12_io_y_sr; // @[package.scala 236:25]
  wire  ppn_data_barrier_12_io_y_pw; // @[package.scala 236:25]
  wire  ppn_data_barrier_12_io_y_px; // @[package.scala 236:25]
  wire  ppn_data_barrier_12_io_y_pr; // @[package.scala 236:25]
  wire  ppn_data_barrier_12_io_y_ppp; // @[package.scala 236:25]
  wire  ppn_data_barrier_12_io_y_pal; // @[package.scala 236:25]
  wire  ppn_data_barrier_12_io_y_paa; // @[package.scala 236:25]
  wire  ppn_data_barrier_12_io_y_eff; // @[package.scala 236:25]
  wire  ppn_data_barrier_12_io_y_c; // @[package.scala 236:25]
  wire [19:0] entries_barrier_io_x_ppn; // @[package.scala 236:25]
  wire  entries_barrier_io_x_u; // @[package.scala 236:25]
  wire  entries_barrier_io_x_ae; // @[package.scala 236:25]
  wire  entries_barrier_io_x_sw; // @[package.scala 236:25]
  wire  entries_barrier_io_x_sx; // @[package.scala 236:25]
  wire  entries_barrier_io_x_sr; // @[package.scala 236:25]
  wire  entries_barrier_io_x_pw; // @[package.scala 236:25]
  wire  entries_barrier_io_x_px; // @[package.scala 236:25]
  wire  entries_barrier_io_x_pr; // @[package.scala 236:25]
  wire  entries_barrier_io_x_ppp; // @[package.scala 236:25]
  wire  entries_barrier_io_x_pal; // @[package.scala 236:25]
  wire  entries_barrier_io_x_paa; // @[package.scala 236:25]
  wire  entries_barrier_io_x_eff; // @[package.scala 236:25]
  wire  entries_barrier_io_x_c; // @[package.scala 236:25]
  wire [19:0] entries_barrier_io_y_ppn; // @[package.scala 236:25]
  wire  entries_barrier_io_y_u; // @[package.scala 236:25]
  wire  entries_barrier_io_y_ae; // @[package.scala 236:25]
  wire  entries_barrier_io_y_sw; // @[package.scala 236:25]
  wire  entries_barrier_io_y_sx; // @[package.scala 236:25]
  wire  entries_barrier_io_y_sr; // @[package.scala 236:25]
  wire  entries_barrier_io_y_pw; // @[package.scala 236:25]
  wire  entries_barrier_io_y_px; // @[package.scala 236:25]
  wire  entries_barrier_io_y_pr; // @[package.scala 236:25]
  wire  entries_barrier_io_y_ppp; // @[package.scala 236:25]
  wire  entries_barrier_io_y_pal; // @[package.scala 236:25]
  wire  entries_barrier_io_y_paa; // @[package.scala 236:25]
  wire  entries_barrier_io_y_eff; // @[package.scala 236:25]
  wire  entries_barrier_io_y_c; // @[package.scala 236:25]
  wire [19:0] entries_barrier_1_io_x_ppn; // @[package.scala 236:25]
  wire  entries_barrier_1_io_x_u; // @[package.scala 236:25]
  wire  entries_barrier_1_io_x_ae; // @[package.scala 236:25]
  wire  entries_barrier_1_io_x_sw; // @[package.scala 236:25]
  wire  entries_barrier_1_io_x_sx; // @[package.scala 236:25]
  wire  entries_barrier_1_io_x_sr; // @[package.scala 236:25]
  wire  entries_barrier_1_io_x_pw; // @[package.scala 236:25]
  wire  entries_barrier_1_io_x_px; // @[package.scala 236:25]
  wire  entries_barrier_1_io_x_pr; // @[package.scala 236:25]
  wire  entries_barrier_1_io_x_ppp; // @[package.scala 236:25]
  wire  entries_barrier_1_io_x_pal; // @[package.scala 236:25]
  wire  entries_barrier_1_io_x_paa; // @[package.scala 236:25]
  wire  entries_barrier_1_io_x_eff; // @[package.scala 236:25]
  wire  entries_barrier_1_io_x_c; // @[package.scala 236:25]
  wire [19:0] entries_barrier_1_io_y_ppn; // @[package.scala 236:25]
  wire  entries_barrier_1_io_y_u; // @[package.scala 236:25]
  wire  entries_barrier_1_io_y_ae; // @[package.scala 236:25]
  wire  entries_barrier_1_io_y_sw; // @[package.scala 236:25]
  wire  entries_barrier_1_io_y_sx; // @[package.scala 236:25]
  wire  entries_barrier_1_io_y_sr; // @[package.scala 236:25]
  wire  entries_barrier_1_io_y_pw; // @[package.scala 236:25]
  wire  entries_barrier_1_io_y_px; // @[package.scala 236:25]
  wire  entries_barrier_1_io_y_pr; // @[package.scala 236:25]
  wire  entries_barrier_1_io_y_ppp; // @[package.scala 236:25]
  wire  entries_barrier_1_io_y_pal; // @[package.scala 236:25]
  wire  entries_barrier_1_io_y_paa; // @[package.scala 236:25]
  wire  entries_barrier_1_io_y_eff; // @[package.scala 236:25]
  wire  entries_barrier_1_io_y_c; // @[package.scala 236:25]
  wire [19:0] entries_barrier_2_io_x_ppn; // @[package.scala 236:25]
  wire  entries_barrier_2_io_x_u; // @[package.scala 236:25]
  wire  entries_barrier_2_io_x_ae; // @[package.scala 236:25]
  wire  entries_barrier_2_io_x_sw; // @[package.scala 236:25]
  wire  entries_barrier_2_io_x_sx; // @[package.scala 236:25]
  wire  entries_barrier_2_io_x_sr; // @[package.scala 236:25]
  wire  entries_barrier_2_io_x_pw; // @[package.scala 236:25]
  wire  entries_barrier_2_io_x_px; // @[package.scala 236:25]
  wire  entries_barrier_2_io_x_pr; // @[package.scala 236:25]
  wire  entries_barrier_2_io_x_ppp; // @[package.scala 236:25]
  wire  entries_barrier_2_io_x_pal; // @[package.scala 236:25]
  wire  entries_barrier_2_io_x_paa; // @[package.scala 236:25]
  wire  entries_barrier_2_io_x_eff; // @[package.scala 236:25]
  wire  entries_barrier_2_io_x_c; // @[package.scala 236:25]
  wire [19:0] entries_barrier_2_io_y_ppn; // @[package.scala 236:25]
  wire  entries_barrier_2_io_y_u; // @[package.scala 236:25]
  wire  entries_barrier_2_io_y_ae; // @[package.scala 236:25]
  wire  entries_barrier_2_io_y_sw; // @[package.scala 236:25]
  wire  entries_barrier_2_io_y_sx; // @[package.scala 236:25]
  wire  entries_barrier_2_io_y_sr; // @[package.scala 236:25]
  wire  entries_barrier_2_io_y_pw; // @[package.scala 236:25]
  wire  entries_barrier_2_io_y_px; // @[package.scala 236:25]
  wire  entries_barrier_2_io_y_pr; // @[package.scala 236:25]
  wire  entries_barrier_2_io_y_ppp; // @[package.scala 236:25]
  wire  entries_barrier_2_io_y_pal; // @[package.scala 236:25]
  wire  entries_barrier_2_io_y_paa; // @[package.scala 236:25]
  wire  entries_barrier_2_io_y_eff; // @[package.scala 236:25]
  wire  entries_barrier_2_io_y_c; // @[package.scala 236:25]
  wire [19:0] entries_barrier_3_io_x_ppn; // @[package.scala 236:25]
  wire  entries_barrier_3_io_x_u; // @[package.scala 236:25]
  wire  entries_barrier_3_io_x_ae; // @[package.scala 236:25]
  wire  entries_barrier_3_io_x_sw; // @[package.scala 236:25]
  wire  entries_barrier_3_io_x_sx; // @[package.scala 236:25]
  wire  entries_barrier_3_io_x_sr; // @[package.scala 236:25]
  wire  entries_barrier_3_io_x_pw; // @[package.scala 236:25]
  wire  entries_barrier_3_io_x_px; // @[package.scala 236:25]
  wire  entries_barrier_3_io_x_pr; // @[package.scala 236:25]
  wire  entries_barrier_3_io_x_ppp; // @[package.scala 236:25]
  wire  entries_barrier_3_io_x_pal; // @[package.scala 236:25]
  wire  entries_barrier_3_io_x_paa; // @[package.scala 236:25]
  wire  entries_barrier_3_io_x_eff; // @[package.scala 236:25]
  wire  entries_barrier_3_io_x_c; // @[package.scala 236:25]
  wire [19:0] entries_barrier_3_io_y_ppn; // @[package.scala 236:25]
  wire  entries_barrier_3_io_y_u; // @[package.scala 236:25]
  wire  entries_barrier_3_io_y_ae; // @[package.scala 236:25]
  wire  entries_barrier_3_io_y_sw; // @[package.scala 236:25]
  wire  entries_barrier_3_io_y_sx; // @[package.scala 236:25]
  wire  entries_barrier_3_io_y_sr; // @[package.scala 236:25]
  wire  entries_barrier_3_io_y_pw; // @[package.scala 236:25]
  wire  entries_barrier_3_io_y_px; // @[package.scala 236:25]
  wire  entries_barrier_3_io_y_pr; // @[package.scala 236:25]
  wire  entries_barrier_3_io_y_ppp; // @[package.scala 236:25]
  wire  entries_barrier_3_io_y_pal; // @[package.scala 236:25]
  wire  entries_barrier_3_io_y_paa; // @[package.scala 236:25]
  wire  entries_barrier_3_io_y_eff; // @[package.scala 236:25]
  wire  entries_barrier_3_io_y_c; // @[package.scala 236:25]
  wire [19:0] entries_barrier_4_io_x_ppn; // @[package.scala 236:25]
  wire  entries_barrier_4_io_x_u; // @[package.scala 236:25]
  wire  entries_barrier_4_io_x_ae; // @[package.scala 236:25]
  wire  entries_barrier_4_io_x_sw; // @[package.scala 236:25]
  wire  entries_barrier_4_io_x_sx; // @[package.scala 236:25]
  wire  entries_barrier_4_io_x_sr; // @[package.scala 236:25]
  wire  entries_barrier_4_io_x_pw; // @[package.scala 236:25]
  wire  entries_barrier_4_io_x_px; // @[package.scala 236:25]
  wire  entries_barrier_4_io_x_pr; // @[package.scala 236:25]
  wire  entries_barrier_4_io_x_ppp; // @[package.scala 236:25]
  wire  entries_barrier_4_io_x_pal; // @[package.scala 236:25]
  wire  entries_barrier_4_io_x_paa; // @[package.scala 236:25]
  wire  entries_barrier_4_io_x_eff; // @[package.scala 236:25]
  wire  entries_barrier_4_io_x_c; // @[package.scala 236:25]
  wire [19:0] entries_barrier_4_io_y_ppn; // @[package.scala 236:25]
  wire  entries_barrier_4_io_y_u; // @[package.scala 236:25]
  wire  entries_barrier_4_io_y_ae; // @[package.scala 236:25]
  wire  entries_barrier_4_io_y_sw; // @[package.scala 236:25]
  wire  entries_barrier_4_io_y_sx; // @[package.scala 236:25]
  wire  entries_barrier_4_io_y_sr; // @[package.scala 236:25]
  wire  entries_barrier_4_io_y_pw; // @[package.scala 236:25]
  wire  entries_barrier_4_io_y_px; // @[package.scala 236:25]
  wire  entries_barrier_4_io_y_pr; // @[package.scala 236:25]
  wire  entries_barrier_4_io_y_ppp; // @[package.scala 236:25]
  wire  entries_barrier_4_io_y_pal; // @[package.scala 236:25]
  wire  entries_barrier_4_io_y_paa; // @[package.scala 236:25]
  wire  entries_barrier_4_io_y_eff; // @[package.scala 236:25]
  wire  entries_barrier_4_io_y_c; // @[package.scala 236:25]
  wire [19:0] entries_barrier_5_io_x_ppn; // @[package.scala 236:25]
  wire  entries_barrier_5_io_x_u; // @[package.scala 236:25]
  wire  entries_barrier_5_io_x_ae; // @[package.scala 236:25]
  wire  entries_barrier_5_io_x_sw; // @[package.scala 236:25]
  wire  entries_barrier_5_io_x_sx; // @[package.scala 236:25]
  wire  entries_barrier_5_io_x_sr; // @[package.scala 236:25]
  wire  entries_barrier_5_io_x_pw; // @[package.scala 236:25]
  wire  entries_barrier_5_io_x_px; // @[package.scala 236:25]
  wire  entries_barrier_5_io_x_pr; // @[package.scala 236:25]
  wire  entries_barrier_5_io_x_ppp; // @[package.scala 236:25]
  wire  entries_barrier_5_io_x_pal; // @[package.scala 236:25]
  wire  entries_barrier_5_io_x_paa; // @[package.scala 236:25]
  wire  entries_barrier_5_io_x_eff; // @[package.scala 236:25]
  wire  entries_barrier_5_io_x_c; // @[package.scala 236:25]
  wire [19:0] entries_barrier_5_io_y_ppn; // @[package.scala 236:25]
  wire  entries_barrier_5_io_y_u; // @[package.scala 236:25]
  wire  entries_barrier_5_io_y_ae; // @[package.scala 236:25]
  wire  entries_barrier_5_io_y_sw; // @[package.scala 236:25]
  wire  entries_barrier_5_io_y_sx; // @[package.scala 236:25]
  wire  entries_barrier_5_io_y_sr; // @[package.scala 236:25]
  wire  entries_barrier_5_io_y_pw; // @[package.scala 236:25]
  wire  entries_barrier_5_io_y_px; // @[package.scala 236:25]
  wire  entries_barrier_5_io_y_pr; // @[package.scala 236:25]
  wire  entries_barrier_5_io_y_ppp; // @[package.scala 236:25]
  wire  entries_barrier_5_io_y_pal; // @[package.scala 236:25]
  wire  entries_barrier_5_io_y_paa; // @[package.scala 236:25]
  wire  entries_barrier_5_io_y_eff; // @[package.scala 236:25]
  wire  entries_barrier_5_io_y_c; // @[package.scala 236:25]
  wire [19:0] entries_barrier_6_io_x_ppn; // @[package.scala 236:25]
  wire  entries_barrier_6_io_x_u; // @[package.scala 236:25]
  wire  entries_barrier_6_io_x_ae; // @[package.scala 236:25]
  wire  entries_barrier_6_io_x_sw; // @[package.scala 236:25]
  wire  entries_barrier_6_io_x_sx; // @[package.scala 236:25]
  wire  entries_barrier_6_io_x_sr; // @[package.scala 236:25]
  wire  entries_barrier_6_io_x_pw; // @[package.scala 236:25]
  wire  entries_barrier_6_io_x_px; // @[package.scala 236:25]
  wire  entries_barrier_6_io_x_pr; // @[package.scala 236:25]
  wire  entries_barrier_6_io_x_ppp; // @[package.scala 236:25]
  wire  entries_barrier_6_io_x_pal; // @[package.scala 236:25]
  wire  entries_barrier_6_io_x_paa; // @[package.scala 236:25]
  wire  entries_barrier_6_io_x_eff; // @[package.scala 236:25]
  wire  entries_barrier_6_io_x_c; // @[package.scala 236:25]
  wire [19:0] entries_barrier_6_io_y_ppn; // @[package.scala 236:25]
  wire  entries_barrier_6_io_y_u; // @[package.scala 236:25]
  wire  entries_barrier_6_io_y_ae; // @[package.scala 236:25]
  wire  entries_barrier_6_io_y_sw; // @[package.scala 236:25]
  wire  entries_barrier_6_io_y_sx; // @[package.scala 236:25]
  wire  entries_barrier_6_io_y_sr; // @[package.scala 236:25]
  wire  entries_barrier_6_io_y_pw; // @[package.scala 236:25]
  wire  entries_barrier_6_io_y_px; // @[package.scala 236:25]
  wire  entries_barrier_6_io_y_pr; // @[package.scala 236:25]
  wire  entries_barrier_6_io_y_ppp; // @[package.scala 236:25]
  wire  entries_barrier_6_io_y_pal; // @[package.scala 236:25]
  wire  entries_barrier_6_io_y_paa; // @[package.scala 236:25]
  wire  entries_barrier_6_io_y_eff; // @[package.scala 236:25]
  wire  entries_barrier_6_io_y_c; // @[package.scala 236:25]
  wire [19:0] entries_barrier_7_io_x_ppn; // @[package.scala 236:25]
  wire  entries_barrier_7_io_x_u; // @[package.scala 236:25]
  wire  entries_barrier_7_io_x_ae; // @[package.scala 236:25]
  wire  entries_barrier_7_io_x_sw; // @[package.scala 236:25]
  wire  entries_barrier_7_io_x_sx; // @[package.scala 236:25]
  wire  entries_barrier_7_io_x_sr; // @[package.scala 236:25]
  wire  entries_barrier_7_io_x_pw; // @[package.scala 236:25]
  wire  entries_barrier_7_io_x_px; // @[package.scala 236:25]
  wire  entries_barrier_7_io_x_pr; // @[package.scala 236:25]
  wire  entries_barrier_7_io_x_ppp; // @[package.scala 236:25]
  wire  entries_barrier_7_io_x_pal; // @[package.scala 236:25]
  wire  entries_barrier_7_io_x_paa; // @[package.scala 236:25]
  wire  entries_barrier_7_io_x_eff; // @[package.scala 236:25]
  wire  entries_barrier_7_io_x_c; // @[package.scala 236:25]
  wire [19:0] entries_barrier_7_io_y_ppn; // @[package.scala 236:25]
  wire  entries_barrier_7_io_y_u; // @[package.scala 236:25]
  wire  entries_barrier_7_io_y_ae; // @[package.scala 236:25]
  wire  entries_barrier_7_io_y_sw; // @[package.scala 236:25]
  wire  entries_barrier_7_io_y_sx; // @[package.scala 236:25]
  wire  entries_barrier_7_io_y_sr; // @[package.scala 236:25]
  wire  entries_barrier_7_io_y_pw; // @[package.scala 236:25]
  wire  entries_barrier_7_io_y_px; // @[package.scala 236:25]
  wire  entries_barrier_7_io_y_pr; // @[package.scala 236:25]
  wire  entries_barrier_7_io_y_ppp; // @[package.scala 236:25]
  wire  entries_barrier_7_io_y_pal; // @[package.scala 236:25]
  wire  entries_barrier_7_io_y_paa; // @[package.scala 236:25]
  wire  entries_barrier_7_io_y_eff; // @[package.scala 236:25]
  wire  entries_barrier_7_io_y_c; // @[package.scala 236:25]
  wire [19:0] entries_barrier_8_io_x_ppn; // @[package.scala 236:25]
  wire  entries_barrier_8_io_x_u; // @[package.scala 236:25]
  wire  entries_barrier_8_io_x_ae; // @[package.scala 236:25]
  wire  entries_barrier_8_io_x_sw; // @[package.scala 236:25]
  wire  entries_barrier_8_io_x_sx; // @[package.scala 236:25]
  wire  entries_barrier_8_io_x_sr; // @[package.scala 236:25]
  wire  entries_barrier_8_io_x_pw; // @[package.scala 236:25]
  wire  entries_barrier_8_io_x_px; // @[package.scala 236:25]
  wire  entries_barrier_8_io_x_pr; // @[package.scala 236:25]
  wire  entries_barrier_8_io_x_ppp; // @[package.scala 236:25]
  wire  entries_barrier_8_io_x_pal; // @[package.scala 236:25]
  wire  entries_barrier_8_io_x_paa; // @[package.scala 236:25]
  wire  entries_barrier_8_io_x_eff; // @[package.scala 236:25]
  wire  entries_barrier_8_io_x_c; // @[package.scala 236:25]
  wire [19:0] entries_barrier_8_io_y_ppn; // @[package.scala 236:25]
  wire  entries_barrier_8_io_y_u; // @[package.scala 236:25]
  wire  entries_barrier_8_io_y_ae; // @[package.scala 236:25]
  wire  entries_barrier_8_io_y_sw; // @[package.scala 236:25]
  wire  entries_barrier_8_io_y_sx; // @[package.scala 236:25]
  wire  entries_barrier_8_io_y_sr; // @[package.scala 236:25]
  wire  entries_barrier_8_io_y_pw; // @[package.scala 236:25]
  wire  entries_barrier_8_io_y_px; // @[package.scala 236:25]
  wire  entries_barrier_8_io_y_pr; // @[package.scala 236:25]
  wire  entries_barrier_8_io_y_ppp; // @[package.scala 236:25]
  wire  entries_barrier_8_io_y_pal; // @[package.scala 236:25]
  wire  entries_barrier_8_io_y_paa; // @[package.scala 236:25]
  wire  entries_barrier_8_io_y_eff; // @[package.scala 236:25]
  wire  entries_barrier_8_io_y_c; // @[package.scala 236:25]
  wire [19:0] entries_barrier_9_io_x_ppn; // @[package.scala 236:25]
  wire  entries_barrier_9_io_x_u; // @[package.scala 236:25]
  wire  entries_barrier_9_io_x_ae; // @[package.scala 236:25]
  wire  entries_barrier_9_io_x_sw; // @[package.scala 236:25]
  wire  entries_barrier_9_io_x_sx; // @[package.scala 236:25]
  wire  entries_barrier_9_io_x_sr; // @[package.scala 236:25]
  wire  entries_barrier_9_io_x_pw; // @[package.scala 236:25]
  wire  entries_barrier_9_io_x_px; // @[package.scala 236:25]
  wire  entries_barrier_9_io_x_pr; // @[package.scala 236:25]
  wire  entries_barrier_9_io_x_ppp; // @[package.scala 236:25]
  wire  entries_barrier_9_io_x_pal; // @[package.scala 236:25]
  wire  entries_barrier_9_io_x_paa; // @[package.scala 236:25]
  wire  entries_barrier_9_io_x_eff; // @[package.scala 236:25]
  wire  entries_barrier_9_io_x_c; // @[package.scala 236:25]
  wire [19:0] entries_barrier_9_io_y_ppn; // @[package.scala 236:25]
  wire  entries_barrier_9_io_y_u; // @[package.scala 236:25]
  wire  entries_barrier_9_io_y_ae; // @[package.scala 236:25]
  wire  entries_barrier_9_io_y_sw; // @[package.scala 236:25]
  wire  entries_barrier_9_io_y_sx; // @[package.scala 236:25]
  wire  entries_barrier_9_io_y_sr; // @[package.scala 236:25]
  wire  entries_barrier_9_io_y_pw; // @[package.scala 236:25]
  wire  entries_barrier_9_io_y_px; // @[package.scala 236:25]
  wire  entries_barrier_9_io_y_pr; // @[package.scala 236:25]
  wire  entries_barrier_9_io_y_ppp; // @[package.scala 236:25]
  wire  entries_barrier_9_io_y_pal; // @[package.scala 236:25]
  wire  entries_barrier_9_io_y_paa; // @[package.scala 236:25]
  wire  entries_barrier_9_io_y_eff; // @[package.scala 236:25]
  wire  entries_barrier_9_io_y_c; // @[package.scala 236:25]
  wire [19:0] entries_barrier_10_io_x_ppn; // @[package.scala 236:25]
  wire  entries_barrier_10_io_x_u; // @[package.scala 236:25]
  wire  entries_barrier_10_io_x_ae; // @[package.scala 236:25]
  wire  entries_barrier_10_io_x_sw; // @[package.scala 236:25]
  wire  entries_barrier_10_io_x_sx; // @[package.scala 236:25]
  wire  entries_barrier_10_io_x_sr; // @[package.scala 236:25]
  wire  entries_barrier_10_io_x_pw; // @[package.scala 236:25]
  wire  entries_barrier_10_io_x_px; // @[package.scala 236:25]
  wire  entries_barrier_10_io_x_pr; // @[package.scala 236:25]
  wire  entries_barrier_10_io_x_ppp; // @[package.scala 236:25]
  wire  entries_barrier_10_io_x_pal; // @[package.scala 236:25]
  wire  entries_barrier_10_io_x_paa; // @[package.scala 236:25]
  wire  entries_barrier_10_io_x_eff; // @[package.scala 236:25]
  wire  entries_barrier_10_io_x_c; // @[package.scala 236:25]
  wire [19:0] entries_barrier_10_io_y_ppn; // @[package.scala 236:25]
  wire  entries_barrier_10_io_y_u; // @[package.scala 236:25]
  wire  entries_barrier_10_io_y_ae; // @[package.scala 236:25]
  wire  entries_barrier_10_io_y_sw; // @[package.scala 236:25]
  wire  entries_barrier_10_io_y_sx; // @[package.scala 236:25]
  wire  entries_barrier_10_io_y_sr; // @[package.scala 236:25]
  wire  entries_barrier_10_io_y_pw; // @[package.scala 236:25]
  wire  entries_barrier_10_io_y_px; // @[package.scala 236:25]
  wire  entries_barrier_10_io_y_pr; // @[package.scala 236:25]
  wire  entries_barrier_10_io_y_ppp; // @[package.scala 236:25]
  wire  entries_barrier_10_io_y_pal; // @[package.scala 236:25]
  wire  entries_barrier_10_io_y_paa; // @[package.scala 236:25]
  wire  entries_barrier_10_io_y_eff; // @[package.scala 236:25]
  wire  entries_barrier_10_io_y_c; // @[package.scala 236:25]
  wire [19:0] entries_barrier_11_io_x_ppn; // @[package.scala 236:25]
  wire  entries_barrier_11_io_x_u; // @[package.scala 236:25]
  wire  entries_barrier_11_io_x_ae; // @[package.scala 236:25]
  wire  entries_barrier_11_io_x_sw; // @[package.scala 236:25]
  wire  entries_barrier_11_io_x_sx; // @[package.scala 236:25]
  wire  entries_barrier_11_io_x_sr; // @[package.scala 236:25]
  wire  entries_barrier_11_io_x_pw; // @[package.scala 236:25]
  wire  entries_barrier_11_io_x_px; // @[package.scala 236:25]
  wire  entries_barrier_11_io_x_pr; // @[package.scala 236:25]
  wire  entries_barrier_11_io_x_ppp; // @[package.scala 236:25]
  wire  entries_barrier_11_io_x_pal; // @[package.scala 236:25]
  wire  entries_barrier_11_io_x_paa; // @[package.scala 236:25]
  wire  entries_barrier_11_io_x_eff; // @[package.scala 236:25]
  wire  entries_barrier_11_io_x_c; // @[package.scala 236:25]
  wire [19:0] entries_barrier_11_io_y_ppn; // @[package.scala 236:25]
  wire  entries_barrier_11_io_y_u; // @[package.scala 236:25]
  wire  entries_barrier_11_io_y_ae; // @[package.scala 236:25]
  wire  entries_barrier_11_io_y_sw; // @[package.scala 236:25]
  wire  entries_barrier_11_io_y_sx; // @[package.scala 236:25]
  wire  entries_barrier_11_io_y_sr; // @[package.scala 236:25]
  wire  entries_barrier_11_io_y_pw; // @[package.scala 236:25]
  wire  entries_barrier_11_io_y_px; // @[package.scala 236:25]
  wire  entries_barrier_11_io_y_pr; // @[package.scala 236:25]
  wire  entries_barrier_11_io_y_ppp; // @[package.scala 236:25]
  wire  entries_barrier_11_io_y_pal; // @[package.scala 236:25]
  wire  entries_barrier_11_io_y_paa; // @[package.scala 236:25]
  wire  entries_barrier_11_io_y_eff; // @[package.scala 236:25]
  wire  entries_barrier_11_io_y_c; // @[package.scala 236:25]
  wire [19:0] entries_barrier_12_io_x_ppn; // @[package.scala 236:25]
  wire  entries_barrier_12_io_x_u; // @[package.scala 236:25]
  wire  entries_barrier_12_io_x_ae; // @[package.scala 236:25]
  wire  entries_barrier_12_io_x_sw; // @[package.scala 236:25]
  wire  entries_barrier_12_io_x_sx; // @[package.scala 236:25]
  wire  entries_barrier_12_io_x_sr; // @[package.scala 236:25]
  wire  entries_barrier_12_io_x_pw; // @[package.scala 236:25]
  wire  entries_barrier_12_io_x_px; // @[package.scala 236:25]
  wire  entries_barrier_12_io_x_pr; // @[package.scala 236:25]
  wire  entries_barrier_12_io_x_ppp; // @[package.scala 236:25]
  wire  entries_barrier_12_io_x_pal; // @[package.scala 236:25]
  wire  entries_barrier_12_io_x_paa; // @[package.scala 236:25]
  wire  entries_barrier_12_io_x_eff; // @[package.scala 236:25]
  wire  entries_barrier_12_io_x_c; // @[package.scala 236:25]
  wire [19:0] entries_barrier_12_io_y_ppn; // @[package.scala 236:25]
  wire  entries_barrier_12_io_y_u; // @[package.scala 236:25]
  wire  entries_barrier_12_io_y_ae; // @[package.scala 236:25]
  wire  entries_barrier_12_io_y_sw; // @[package.scala 236:25]
  wire  entries_barrier_12_io_y_sx; // @[package.scala 236:25]
  wire  entries_barrier_12_io_y_sr; // @[package.scala 236:25]
  wire  entries_barrier_12_io_y_pw; // @[package.scala 236:25]
  wire  entries_barrier_12_io_y_px; // @[package.scala 236:25]
  wire  entries_barrier_12_io_y_pr; // @[package.scala 236:25]
  wire  entries_barrier_12_io_y_ppp; // @[package.scala 236:25]
  wire  entries_barrier_12_io_y_pal; // @[package.scala 236:25]
  wire  entries_barrier_12_io_y_paa; // @[package.scala 236:25]
  wire  entries_barrier_12_io_y_eff; // @[package.scala 236:25]
  wire  entries_barrier_12_io_y_c; // @[package.scala 236:25]
  wire [19:0] normal_entries_barrier_io_x_ppn; // @[package.scala 236:25]
  wire  normal_entries_barrier_io_x_u; // @[package.scala 236:25]
  wire  normal_entries_barrier_io_x_ae; // @[package.scala 236:25]
  wire  normal_entries_barrier_io_x_sw; // @[package.scala 236:25]
  wire  normal_entries_barrier_io_x_sx; // @[package.scala 236:25]
  wire  normal_entries_barrier_io_x_sr; // @[package.scala 236:25]
  wire  normal_entries_barrier_io_x_pw; // @[package.scala 236:25]
  wire  normal_entries_barrier_io_x_px; // @[package.scala 236:25]
  wire  normal_entries_barrier_io_x_pr; // @[package.scala 236:25]
  wire  normal_entries_barrier_io_x_ppp; // @[package.scala 236:25]
  wire  normal_entries_barrier_io_x_pal; // @[package.scala 236:25]
  wire  normal_entries_barrier_io_x_paa; // @[package.scala 236:25]
  wire  normal_entries_barrier_io_x_eff; // @[package.scala 236:25]
  wire  normal_entries_barrier_io_x_c; // @[package.scala 236:25]
  wire [19:0] normal_entries_barrier_io_y_ppn; // @[package.scala 236:25]
  wire  normal_entries_barrier_io_y_u; // @[package.scala 236:25]
  wire  normal_entries_barrier_io_y_ae; // @[package.scala 236:25]
  wire  normal_entries_barrier_io_y_sw; // @[package.scala 236:25]
  wire  normal_entries_barrier_io_y_sx; // @[package.scala 236:25]
  wire  normal_entries_barrier_io_y_sr; // @[package.scala 236:25]
  wire  normal_entries_barrier_io_y_pw; // @[package.scala 236:25]
  wire  normal_entries_barrier_io_y_px; // @[package.scala 236:25]
  wire  normal_entries_barrier_io_y_pr; // @[package.scala 236:25]
  wire  normal_entries_barrier_io_y_ppp; // @[package.scala 236:25]
  wire  normal_entries_barrier_io_y_pal; // @[package.scala 236:25]
  wire  normal_entries_barrier_io_y_paa; // @[package.scala 236:25]
  wire  normal_entries_barrier_io_y_eff; // @[package.scala 236:25]
  wire  normal_entries_barrier_io_y_c; // @[package.scala 236:25]
  wire [19:0] normal_entries_barrier_1_io_x_ppn; // @[package.scala 236:25]
  wire  normal_entries_barrier_1_io_x_u; // @[package.scala 236:25]
  wire  normal_entries_barrier_1_io_x_ae; // @[package.scala 236:25]
  wire  normal_entries_barrier_1_io_x_sw; // @[package.scala 236:25]
  wire  normal_entries_barrier_1_io_x_sx; // @[package.scala 236:25]
  wire  normal_entries_barrier_1_io_x_sr; // @[package.scala 236:25]
  wire  normal_entries_barrier_1_io_x_pw; // @[package.scala 236:25]
  wire  normal_entries_barrier_1_io_x_px; // @[package.scala 236:25]
  wire  normal_entries_barrier_1_io_x_pr; // @[package.scala 236:25]
  wire  normal_entries_barrier_1_io_x_ppp; // @[package.scala 236:25]
  wire  normal_entries_barrier_1_io_x_pal; // @[package.scala 236:25]
  wire  normal_entries_barrier_1_io_x_paa; // @[package.scala 236:25]
  wire  normal_entries_barrier_1_io_x_eff; // @[package.scala 236:25]
  wire  normal_entries_barrier_1_io_x_c; // @[package.scala 236:25]
  wire [19:0] normal_entries_barrier_1_io_y_ppn; // @[package.scala 236:25]
  wire  normal_entries_barrier_1_io_y_u; // @[package.scala 236:25]
  wire  normal_entries_barrier_1_io_y_ae; // @[package.scala 236:25]
  wire  normal_entries_barrier_1_io_y_sw; // @[package.scala 236:25]
  wire  normal_entries_barrier_1_io_y_sx; // @[package.scala 236:25]
  wire  normal_entries_barrier_1_io_y_sr; // @[package.scala 236:25]
  wire  normal_entries_barrier_1_io_y_pw; // @[package.scala 236:25]
  wire  normal_entries_barrier_1_io_y_px; // @[package.scala 236:25]
  wire  normal_entries_barrier_1_io_y_pr; // @[package.scala 236:25]
  wire  normal_entries_barrier_1_io_y_ppp; // @[package.scala 236:25]
  wire  normal_entries_barrier_1_io_y_pal; // @[package.scala 236:25]
  wire  normal_entries_barrier_1_io_y_paa; // @[package.scala 236:25]
  wire  normal_entries_barrier_1_io_y_eff; // @[package.scala 236:25]
  wire  normal_entries_barrier_1_io_y_c; // @[package.scala 236:25]
  wire [19:0] normal_entries_barrier_2_io_x_ppn; // @[package.scala 236:25]
  wire  normal_entries_barrier_2_io_x_u; // @[package.scala 236:25]
  wire  normal_entries_barrier_2_io_x_ae; // @[package.scala 236:25]
  wire  normal_entries_barrier_2_io_x_sw; // @[package.scala 236:25]
  wire  normal_entries_barrier_2_io_x_sx; // @[package.scala 236:25]
  wire  normal_entries_barrier_2_io_x_sr; // @[package.scala 236:25]
  wire  normal_entries_barrier_2_io_x_pw; // @[package.scala 236:25]
  wire  normal_entries_barrier_2_io_x_px; // @[package.scala 236:25]
  wire  normal_entries_barrier_2_io_x_pr; // @[package.scala 236:25]
  wire  normal_entries_barrier_2_io_x_ppp; // @[package.scala 236:25]
  wire  normal_entries_barrier_2_io_x_pal; // @[package.scala 236:25]
  wire  normal_entries_barrier_2_io_x_paa; // @[package.scala 236:25]
  wire  normal_entries_barrier_2_io_x_eff; // @[package.scala 236:25]
  wire  normal_entries_barrier_2_io_x_c; // @[package.scala 236:25]
  wire [19:0] normal_entries_barrier_2_io_y_ppn; // @[package.scala 236:25]
  wire  normal_entries_barrier_2_io_y_u; // @[package.scala 236:25]
  wire  normal_entries_barrier_2_io_y_ae; // @[package.scala 236:25]
  wire  normal_entries_barrier_2_io_y_sw; // @[package.scala 236:25]
  wire  normal_entries_barrier_2_io_y_sx; // @[package.scala 236:25]
  wire  normal_entries_barrier_2_io_y_sr; // @[package.scala 236:25]
  wire  normal_entries_barrier_2_io_y_pw; // @[package.scala 236:25]
  wire  normal_entries_barrier_2_io_y_px; // @[package.scala 236:25]
  wire  normal_entries_barrier_2_io_y_pr; // @[package.scala 236:25]
  wire  normal_entries_barrier_2_io_y_ppp; // @[package.scala 236:25]
  wire  normal_entries_barrier_2_io_y_pal; // @[package.scala 236:25]
  wire  normal_entries_barrier_2_io_y_paa; // @[package.scala 236:25]
  wire  normal_entries_barrier_2_io_y_eff; // @[package.scala 236:25]
  wire  normal_entries_barrier_2_io_y_c; // @[package.scala 236:25]
  wire [19:0] normal_entries_barrier_3_io_x_ppn; // @[package.scala 236:25]
  wire  normal_entries_barrier_3_io_x_u; // @[package.scala 236:25]
  wire  normal_entries_barrier_3_io_x_ae; // @[package.scala 236:25]
  wire  normal_entries_barrier_3_io_x_sw; // @[package.scala 236:25]
  wire  normal_entries_barrier_3_io_x_sx; // @[package.scala 236:25]
  wire  normal_entries_barrier_3_io_x_sr; // @[package.scala 236:25]
  wire  normal_entries_barrier_3_io_x_pw; // @[package.scala 236:25]
  wire  normal_entries_barrier_3_io_x_px; // @[package.scala 236:25]
  wire  normal_entries_barrier_3_io_x_pr; // @[package.scala 236:25]
  wire  normal_entries_barrier_3_io_x_ppp; // @[package.scala 236:25]
  wire  normal_entries_barrier_3_io_x_pal; // @[package.scala 236:25]
  wire  normal_entries_barrier_3_io_x_paa; // @[package.scala 236:25]
  wire  normal_entries_barrier_3_io_x_eff; // @[package.scala 236:25]
  wire  normal_entries_barrier_3_io_x_c; // @[package.scala 236:25]
  wire [19:0] normal_entries_barrier_3_io_y_ppn; // @[package.scala 236:25]
  wire  normal_entries_barrier_3_io_y_u; // @[package.scala 236:25]
  wire  normal_entries_barrier_3_io_y_ae; // @[package.scala 236:25]
  wire  normal_entries_barrier_3_io_y_sw; // @[package.scala 236:25]
  wire  normal_entries_barrier_3_io_y_sx; // @[package.scala 236:25]
  wire  normal_entries_barrier_3_io_y_sr; // @[package.scala 236:25]
  wire  normal_entries_barrier_3_io_y_pw; // @[package.scala 236:25]
  wire  normal_entries_barrier_3_io_y_px; // @[package.scala 236:25]
  wire  normal_entries_barrier_3_io_y_pr; // @[package.scala 236:25]
  wire  normal_entries_barrier_3_io_y_ppp; // @[package.scala 236:25]
  wire  normal_entries_barrier_3_io_y_pal; // @[package.scala 236:25]
  wire  normal_entries_barrier_3_io_y_paa; // @[package.scala 236:25]
  wire  normal_entries_barrier_3_io_y_eff; // @[package.scala 236:25]
  wire  normal_entries_barrier_3_io_y_c; // @[package.scala 236:25]
  wire [19:0] normal_entries_barrier_4_io_x_ppn; // @[package.scala 236:25]
  wire  normal_entries_barrier_4_io_x_u; // @[package.scala 236:25]
  wire  normal_entries_barrier_4_io_x_ae; // @[package.scala 236:25]
  wire  normal_entries_barrier_4_io_x_sw; // @[package.scala 236:25]
  wire  normal_entries_barrier_4_io_x_sx; // @[package.scala 236:25]
  wire  normal_entries_barrier_4_io_x_sr; // @[package.scala 236:25]
  wire  normal_entries_barrier_4_io_x_pw; // @[package.scala 236:25]
  wire  normal_entries_barrier_4_io_x_px; // @[package.scala 236:25]
  wire  normal_entries_barrier_4_io_x_pr; // @[package.scala 236:25]
  wire  normal_entries_barrier_4_io_x_ppp; // @[package.scala 236:25]
  wire  normal_entries_barrier_4_io_x_pal; // @[package.scala 236:25]
  wire  normal_entries_barrier_4_io_x_paa; // @[package.scala 236:25]
  wire  normal_entries_barrier_4_io_x_eff; // @[package.scala 236:25]
  wire  normal_entries_barrier_4_io_x_c; // @[package.scala 236:25]
  wire [19:0] normal_entries_barrier_4_io_y_ppn; // @[package.scala 236:25]
  wire  normal_entries_barrier_4_io_y_u; // @[package.scala 236:25]
  wire  normal_entries_barrier_4_io_y_ae; // @[package.scala 236:25]
  wire  normal_entries_barrier_4_io_y_sw; // @[package.scala 236:25]
  wire  normal_entries_barrier_4_io_y_sx; // @[package.scala 236:25]
  wire  normal_entries_barrier_4_io_y_sr; // @[package.scala 236:25]
  wire  normal_entries_barrier_4_io_y_pw; // @[package.scala 236:25]
  wire  normal_entries_barrier_4_io_y_px; // @[package.scala 236:25]
  wire  normal_entries_barrier_4_io_y_pr; // @[package.scala 236:25]
  wire  normal_entries_barrier_4_io_y_ppp; // @[package.scala 236:25]
  wire  normal_entries_barrier_4_io_y_pal; // @[package.scala 236:25]
  wire  normal_entries_barrier_4_io_y_paa; // @[package.scala 236:25]
  wire  normal_entries_barrier_4_io_y_eff; // @[package.scala 236:25]
  wire  normal_entries_barrier_4_io_y_c; // @[package.scala 236:25]
  wire [19:0] normal_entries_barrier_5_io_x_ppn; // @[package.scala 236:25]
  wire  normal_entries_barrier_5_io_x_u; // @[package.scala 236:25]
  wire  normal_entries_barrier_5_io_x_ae; // @[package.scala 236:25]
  wire  normal_entries_barrier_5_io_x_sw; // @[package.scala 236:25]
  wire  normal_entries_barrier_5_io_x_sx; // @[package.scala 236:25]
  wire  normal_entries_barrier_5_io_x_sr; // @[package.scala 236:25]
  wire  normal_entries_barrier_5_io_x_pw; // @[package.scala 236:25]
  wire  normal_entries_barrier_5_io_x_px; // @[package.scala 236:25]
  wire  normal_entries_barrier_5_io_x_pr; // @[package.scala 236:25]
  wire  normal_entries_barrier_5_io_x_ppp; // @[package.scala 236:25]
  wire  normal_entries_barrier_5_io_x_pal; // @[package.scala 236:25]
  wire  normal_entries_barrier_5_io_x_paa; // @[package.scala 236:25]
  wire  normal_entries_barrier_5_io_x_eff; // @[package.scala 236:25]
  wire  normal_entries_barrier_5_io_x_c; // @[package.scala 236:25]
  wire [19:0] normal_entries_barrier_5_io_y_ppn; // @[package.scala 236:25]
  wire  normal_entries_barrier_5_io_y_u; // @[package.scala 236:25]
  wire  normal_entries_barrier_5_io_y_ae; // @[package.scala 236:25]
  wire  normal_entries_barrier_5_io_y_sw; // @[package.scala 236:25]
  wire  normal_entries_barrier_5_io_y_sx; // @[package.scala 236:25]
  wire  normal_entries_barrier_5_io_y_sr; // @[package.scala 236:25]
  wire  normal_entries_barrier_5_io_y_pw; // @[package.scala 236:25]
  wire  normal_entries_barrier_5_io_y_px; // @[package.scala 236:25]
  wire  normal_entries_barrier_5_io_y_pr; // @[package.scala 236:25]
  wire  normal_entries_barrier_5_io_y_ppp; // @[package.scala 236:25]
  wire  normal_entries_barrier_5_io_y_pal; // @[package.scala 236:25]
  wire  normal_entries_barrier_5_io_y_paa; // @[package.scala 236:25]
  wire  normal_entries_barrier_5_io_y_eff; // @[package.scala 236:25]
  wire  normal_entries_barrier_5_io_y_c; // @[package.scala 236:25]
  wire [19:0] normal_entries_barrier_6_io_x_ppn; // @[package.scala 236:25]
  wire  normal_entries_barrier_6_io_x_u; // @[package.scala 236:25]
  wire  normal_entries_barrier_6_io_x_ae; // @[package.scala 236:25]
  wire  normal_entries_barrier_6_io_x_sw; // @[package.scala 236:25]
  wire  normal_entries_barrier_6_io_x_sx; // @[package.scala 236:25]
  wire  normal_entries_barrier_6_io_x_sr; // @[package.scala 236:25]
  wire  normal_entries_barrier_6_io_x_pw; // @[package.scala 236:25]
  wire  normal_entries_barrier_6_io_x_px; // @[package.scala 236:25]
  wire  normal_entries_barrier_6_io_x_pr; // @[package.scala 236:25]
  wire  normal_entries_barrier_6_io_x_ppp; // @[package.scala 236:25]
  wire  normal_entries_barrier_6_io_x_pal; // @[package.scala 236:25]
  wire  normal_entries_barrier_6_io_x_paa; // @[package.scala 236:25]
  wire  normal_entries_barrier_6_io_x_eff; // @[package.scala 236:25]
  wire  normal_entries_barrier_6_io_x_c; // @[package.scala 236:25]
  wire [19:0] normal_entries_barrier_6_io_y_ppn; // @[package.scala 236:25]
  wire  normal_entries_barrier_6_io_y_u; // @[package.scala 236:25]
  wire  normal_entries_barrier_6_io_y_ae; // @[package.scala 236:25]
  wire  normal_entries_barrier_6_io_y_sw; // @[package.scala 236:25]
  wire  normal_entries_barrier_6_io_y_sx; // @[package.scala 236:25]
  wire  normal_entries_barrier_6_io_y_sr; // @[package.scala 236:25]
  wire  normal_entries_barrier_6_io_y_pw; // @[package.scala 236:25]
  wire  normal_entries_barrier_6_io_y_px; // @[package.scala 236:25]
  wire  normal_entries_barrier_6_io_y_pr; // @[package.scala 236:25]
  wire  normal_entries_barrier_6_io_y_ppp; // @[package.scala 236:25]
  wire  normal_entries_barrier_6_io_y_pal; // @[package.scala 236:25]
  wire  normal_entries_barrier_6_io_y_paa; // @[package.scala 236:25]
  wire  normal_entries_barrier_6_io_y_eff; // @[package.scala 236:25]
  wire  normal_entries_barrier_6_io_y_c; // @[package.scala 236:25]
  wire [19:0] normal_entries_barrier_7_io_x_ppn; // @[package.scala 236:25]
  wire  normal_entries_barrier_7_io_x_u; // @[package.scala 236:25]
  wire  normal_entries_barrier_7_io_x_ae; // @[package.scala 236:25]
  wire  normal_entries_barrier_7_io_x_sw; // @[package.scala 236:25]
  wire  normal_entries_barrier_7_io_x_sx; // @[package.scala 236:25]
  wire  normal_entries_barrier_7_io_x_sr; // @[package.scala 236:25]
  wire  normal_entries_barrier_7_io_x_pw; // @[package.scala 236:25]
  wire  normal_entries_barrier_7_io_x_px; // @[package.scala 236:25]
  wire  normal_entries_barrier_7_io_x_pr; // @[package.scala 236:25]
  wire  normal_entries_barrier_7_io_x_ppp; // @[package.scala 236:25]
  wire  normal_entries_barrier_7_io_x_pal; // @[package.scala 236:25]
  wire  normal_entries_barrier_7_io_x_paa; // @[package.scala 236:25]
  wire  normal_entries_barrier_7_io_x_eff; // @[package.scala 236:25]
  wire  normal_entries_barrier_7_io_x_c; // @[package.scala 236:25]
  wire [19:0] normal_entries_barrier_7_io_y_ppn; // @[package.scala 236:25]
  wire  normal_entries_barrier_7_io_y_u; // @[package.scala 236:25]
  wire  normal_entries_barrier_7_io_y_ae; // @[package.scala 236:25]
  wire  normal_entries_barrier_7_io_y_sw; // @[package.scala 236:25]
  wire  normal_entries_barrier_7_io_y_sx; // @[package.scala 236:25]
  wire  normal_entries_barrier_7_io_y_sr; // @[package.scala 236:25]
  wire  normal_entries_barrier_7_io_y_pw; // @[package.scala 236:25]
  wire  normal_entries_barrier_7_io_y_px; // @[package.scala 236:25]
  wire  normal_entries_barrier_7_io_y_pr; // @[package.scala 236:25]
  wire  normal_entries_barrier_7_io_y_ppp; // @[package.scala 236:25]
  wire  normal_entries_barrier_7_io_y_pal; // @[package.scala 236:25]
  wire  normal_entries_barrier_7_io_y_paa; // @[package.scala 236:25]
  wire  normal_entries_barrier_7_io_y_eff; // @[package.scala 236:25]
  wire  normal_entries_barrier_7_io_y_c; // @[package.scala 236:25]
  wire [19:0] normal_entries_barrier_8_io_x_ppn; // @[package.scala 236:25]
  wire  normal_entries_barrier_8_io_x_u; // @[package.scala 236:25]
  wire  normal_entries_barrier_8_io_x_ae; // @[package.scala 236:25]
  wire  normal_entries_barrier_8_io_x_sw; // @[package.scala 236:25]
  wire  normal_entries_barrier_8_io_x_sx; // @[package.scala 236:25]
  wire  normal_entries_barrier_8_io_x_sr; // @[package.scala 236:25]
  wire  normal_entries_barrier_8_io_x_pw; // @[package.scala 236:25]
  wire  normal_entries_barrier_8_io_x_px; // @[package.scala 236:25]
  wire  normal_entries_barrier_8_io_x_pr; // @[package.scala 236:25]
  wire  normal_entries_barrier_8_io_x_ppp; // @[package.scala 236:25]
  wire  normal_entries_barrier_8_io_x_pal; // @[package.scala 236:25]
  wire  normal_entries_barrier_8_io_x_paa; // @[package.scala 236:25]
  wire  normal_entries_barrier_8_io_x_eff; // @[package.scala 236:25]
  wire  normal_entries_barrier_8_io_x_c; // @[package.scala 236:25]
  wire [19:0] normal_entries_barrier_8_io_y_ppn; // @[package.scala 236:25]
  wire  normal_entries_barrier_8_io_y_u; // @[package.scala 236:25]
  wire  normal_entries_barrier_8_io_y_ae; // @[package.scala 236:25]
  wire  normal_entries_barrier_8_io_y_sw; // @[package.scala 236:25]
  wire  normal_entries_barrier_8_io_y_sx; // @[package.scala 236:25]
  wire  normal_entries_barrier_8_io_y_sr; // @[package.scala 236:25]
  wire  normal_entries_barrier_8_io_y_pw; // @[package.scala 236:25]
  wire  normal_entries_barrier_8_io_y_px; // @[package.scala 236:25]
  wire  normal_entries_barrier_8_io_y_pr; // @[package.scala 236:25]
  wire  normal_entries_barrier_8_io_y_ppp; // @[package.scala 236:25]
  wire  normal_entries_barrier_8_io_y_pal; // @[package.scala 236:25]
  wire  normal_entries_barrier_8_io_y_paa; // @[package.scala 236:25]
  wire  normal_entries_barrier_8_io_y_eff; // @[package.scala 236:25]
  wire  normal_entries_barrier_8_io_y_c; // @[package.scala 236:25]
  wire [19:0] normal_entries_barrier_9_io_x_ppn; // @[package.scala 236:25]
  wire  normal_entries_barrier_9_io_x_u; // @[package.scala 236:25]
  wire  normal_entries_barrier_9_io_x_ae; // @[package.scala 236:25]
  wire  normal_entries_barrier_9_io_x_sw; // @[package.scala 236:25]
  wire  normal_entries_barrier_9_io_x_sx; // @[package.scala 236:25]
  wire  normal_entries_barrier_9_io_x_sr; // @[package.scala 236:25]
  wire  normal_entries_barrier_9_io_x_pw; // @[package.scala 236:25]
  wire  normal_entries_barrier_9_io_x_px; // @[package.scala 236:25]
  wire  normal_entries_barrier_9_io_x_pr; // @[package.scala 236:25]
  wire  normal_entries_barrier_9_io_x_ppp; // @[package.scala 236:25]
  wire  normal_entries_barrier_9_io_x_pal; // @[package.scala 236:25]
  wire  normal_entries_barrier_9_io_x_paa; // @[package.scala 236:25]
  wire  normal_entries_barrier_9_io_x_eff; // @[package.scala 236:25]
  wire  normal_entries_barrier_9_io_x_c; // @[package.scala 236:25]
  wire [19:0] normal_entries_barrier_9_io_y_ppn; // @[package.scala 236:25]
  wire  normal_entries_barrier_9_io_y_u; // @[package.scala 236:25]
  wire  normal_entries_barrier_9_io_y_ae; // @[package.scala 236:25]
  wire  normal_entries_barrier_9_io_y_sw; // @[package.scala 236:25]
  wire  normal_entries_barrier_9_io_y_sx; // @[package.scala 236:25]
  wire  normal_entries_barrier_9_io_y_sr; // @[package.scala 236:25]
  wire  normal_entries_barrier_9_io_y_pw; // @[package.scala 236:25]
  wire  normal_entries_barrier_9_io_y_px; // @[package.scala 236:25]
  wire  normal_entries_barrier_9_io_y_pr; // @[package.scala 236:25]
  wire  normal_entries_barrier_9_io_y_ppp; // @[package.scala 236:25]
  wire  normal_entries_barrier_9_io_y_pal; // @[package.scala 236:25]
  wire  normal_entries_barrier_9_io_y_paa; // @[package.scala 236:25]
  wire  normal_entries_barrier_9_io_y_eff; // @[package.scala 236:25]
  wire  normal_entries_barrier_9_io_y_c; // @[package.scala 236:25]
  wire [19:0] normal_entries_barrier_10_io_x_ppn; // @[package.scala 236:25]
  wire  normal_entries_barrier_10_io_x_u; // @[package.scala 236:25]
  wire  normal_entries_barrier_10_io_x_ae; // @[package.scala 236:25]
  wire  normal_entries_barrier_10_io_x_sw; // @[package.scala 236:25]
  wire  normal_entries_barrier_10_io_x_sx; // @[package.scala 236:25]
  wire  normal_entries_barrier_10_io_x_sr; // @[package.scala 236:25]
  wire  normal_entries_barrier_10_io_x_pw; // @[package.scala 236:25]
  wire  normal_entries_barrier_10_io_x_px; // @[package.scala 236:25]
  wire  normal_entries_barrier_10_io_x_pr; // @[package.scala 236:25]
  wire  normal_entries_barrier_10_io_x_ppp; // @[package.scala 236:25]
  wire  normal_entries_barrier_10_io_x_pal; // @[package.scala 236:25]
  wire  normal_entries_barrier_10_io_x_paa; // @[package.scala 236:25]
  wire  normal_entries_barrier_10_io_x_eff; // @[package.scala 236:25]
  wire  normal_entries_barrier_10_io_x_c; // @[package.scala 236:25]
  wire [19:0] normal_entries_barrier_10_io_y_ppn; // @[package.scala 236:25]
  wire  normal_entries_barrier_10_io_y_u; // @[package.scala 236:25]
  wire  normal_entries_barrier_10_io_y_ae; // @[package.scala 236:25]
  wire  normal_entries_barrier_10_io_y_sw; // @[package.scala 236:25]
  wire  normal_entries_barrier_10_io_y_sx; // @[package.scala 236:25]
  wire  normal_entries_barrier_10_io_y_sr; // @[package.scala 236:25]
  wire  normal_entries_barrier_10_io_y_pw; // @[package.scala 236:25]
  wire  normal_entries_barrier_10_io_y_px; // @[package.scala 236:25]
  wire  normal_entries_barrier_10_io_y_pr; // @[package.scala 236:25]
  wire  normal_entries_barrier_10_io_y_ppp; // @[package.scala 236:25]
  wire  normal_entries_barrier_10_io_y_pal; // @[package.scala 236:25]
  wire  normal_entries_barrier_10_io_y_paa; // @[package.scala 236:25]
  wire  normal_entries_barrier_10_io_y_eff; // @[package.scala 236:25]
  wire  normal_entries_barrier_10_io_y_c; // @[package.scala 236:25]
  wire [19:0] normal_entries_barrier_11_io_x_ppn; // @[package.scala 236:25]
  wire  normal_entries_barrier_11_io_x_u; // @[package.scala 236:25]
  wire  normal_entries_barrier_11_io_x_ae; // @[package.scala 236:25]
  wire  normal_entries_barrier_11_io_x_sw; // @[package.scala 236:25]
  wire  normal_entries_barrier_11_io_x_sx; // @[package.scala 236:25]
  wire  normal_entries_barrier_11_io_x_sr; // @[package.scala 236:25]
  wire  normal_entries_barrier_11_io_x_pw; // @[package.scala 236:25]
  wire  normal_entries_barrier_11_io_x_px; // @[package.scala 236:25]
  wire  normal_entries_barrier_11_io_x_pr; // @[package.scala 236:25]
  wire  normal_entries_barrier_11_io_x_ppp; // @[package.scala 236:25]
  wire  normal_entries_barrier_11_io_x_pal; // @[package.scala 236:25]
  wire  normal_entries_barrier_11_io_x_paa; // @[package.scala 236:25]
  wire  normal_entries_barrier_11_io_x_eff; // @[package.scala 236:25]
  wire  normal_entries_barrier_11_io_x_c; // @[package.scala 236:25]
  wire [19:0] normal_entries_barrier_11_io_y_ppn; // @[package.scala 236:25]
  wire  normal_entries_barrier_11_io_y_u; // @[package.scala 236:25]
  wire  normal_entries_barrier_11_io_y_ae; // @[package.scala 236:25]
  wire  normal_entries_barrier_11_io_y_sw; // @[package.scala 236:25]
  wire  normal_entries_barrier_11_io_y_sx; // @[package.scala 236:25]
  wire  normal_entries_barrier_11_io_y_sr; // @[package.scala 236:25]
  wire  normal_entries_barrier_11_io_y_pw; // @[package.scala 236:25]
  wire  normal_entries_barrier_11_io_y_px; // @[package.scala 236:25]
  wire  normal_entries_barrier_11_io_y_pr; // @[package.scala 236:25]
  wire  normal_entries_barrier_11_io_y_ppp; // @[package.scala 236:25]
  wire  normal_entries_barrier_11_io_y_pal; // @[package.scala 236:25]
  wire  normal_entries_barrier_11_io_y_paa; // @[package.scala 236:25]
  wire  normal_entries_barrier_11_io_y_eff; // @[package.scala 236:25]
  wire  normal_entries_barrier_11_io_y_c; // @[package.scala 236:25]
  reg [26:0] sectored_entries_0_tag; // @[TLB.scala 162:29]
  reg [34:0] sectored_entries_0_data_0; // @[TLB.scala 162:29]
  reg [34:0] sectored_entries_0_data_1; // @[TLB.scala 162:29]
  reg [34:0] sectored_entries_0_data_2; // @[TLB.scala 162:29]
  reg [34:0] sectored_entries_0_data_3; // @[TLB.scala 162:29]
  reg  sectored_entries_0_valid_0; // @[TLB.scala 162:29]
  reg  sectored_entries_0_valid_1; // @[TLB.scala 162:29]
  reg  sectored_entries_0_valid_2; // @[TLB.scala 162:29]
  reg  sectored_entries_0_valid_3; // @[TLB.scala 162:29]
  reg [26:0] sectored_entries_1_tag; // @[TLB.scala 162:29]
  reg [34:0] sectored_entries_1_data_0; // @[TLB.scala 162:29]
  reg [34:0] sectored_entries_1_data_1; // @[TLB.scala 162:29]
  reg [34:0] sectored_entries_1_data_2; // @[TLB.scala 162:29]
  reg [34:0] sectored_entries_1_data_3; // @[TLB.scala 162:29]
  reg  sectored_entries_1_valid_0; // @[TLB.scala 162:29]
  reg  sectored_entries_1_valid_1; // @[TLB.scala 162:29]
  reg  sectored_entries_1_valid_2; // @[TLB.scala 162:29]
  reg  sectored_entries_1_valid_3; // @[TLB.scala 162:29]
  reg [26:0] sectored_entries_2_tag; // @[TLB.scala 162:29]
  reg [34:0] sectored_entries_2_data_0; // @[TLB.scala 162:29]
  reg [34:0] sectored_entries_2_data_1; // @[TLB.scala 162:29]
  reg [34:0] sectored_entries_2_data_2; // @[TLB.scala 162:29]
  reg [34:0] sectored_entries_2_data_3; // @[TLB.scala 162:29]
  reg  sectored_entries_2_valid_0; // @[TLB.scala 162:29]
  reg  sectored_entries_2_valid_1; // @[TLB.scala 162:29]
  reg  sectored_entries_2_valid_2; // @[TLB.scala 162:29]
  reg  sectored_entries_2_valid_3; // @[TLB.scala 162:29]
  reg [26:0] sectored_entries_3_tag; // @[TLB.scala 162:29]
  reg [34:0] sectored_entries_3_data_0; // @[TLB.scala 162:29]
  reg [34:0] sectored_entries_3_data_1; // @[TLB.scala 162:29]
  reg [34:0] sectored_entries_3_data_2; // @[TLB.scala 162:29]
  reg [34:0] sectored_entries_3_data_3; // @[TLB.scala 162:29]
  reg  sectored_entries_3_valid_0; // @[TLB.scala 162:29]
  reg  sectored_entries_3_valid_1; // @[TLB.scala 162:29]
  reg  sectored_entries_3_valid_2; // @[TLB.scala 162:29]
  reg  sectored_entries_3_valid_3; // @[TLB.scala 162:29]
  reg [26:0] sectored_entries_4_tag; // @[TLB.scala 162:29]
  reg [34:0] sectored_entries_4_data_0; // @[TLB.scala 162:29]
  reg [34:0] sectored_entries_4_data_1; // @[TLB.scala 162:29]
  reg [34:0] sectored_entries_4_data_2; // @[TLB.scala 162:29]
  reg [34:0] sectored_entries_4_data_3; // @[TLB.scala 162:29]
  reg  sectored_entries_4_valid_0; // @[TLB.scala 162:29]
  reg  sectored_entries_4_valid_1; // @[TLB.scala 162:29]
  reg  sectored_entries_4_valid_2; // @[TLB.scala 162:29]
  reg  sectored_entries_4_valid_3; // @[TLB.scala 162:29]
  reg [26:0] sectored_entries_5_tag; // @[TLB.scala 162:29]
  reg [34:0] sectored_entries_5_data_0; // @[TLB.scala 162:29]
  reg [34:0] sectored_entries_5_data_1; // @[TLB.scala 162:29]
  reg [34:0] sectored_entries_5_data_2; // @[TLB.scala 162:29]
  reg [34:0] sectored_entries_5_data_3; // @[TLB.scala 162:29]
  reg  sectored_entries_5_valid_0; // @[TLB.scala 162:29]
  reg  sectored_entries_5_valid_1; // @[TLB.scala 162:29]
  reg  sectored_entries_5_valid_2; // @[TLB.scala 162:29]
  reg  sectored_entries_5_valid_3; // @[TLB.scala 162:29]
  reg [26:0] sectored_entries_6_tag; // @[TLB.scala 162:29]
  reg [34:0] sectored_entries_6_data_0; // @[TLB.scala 162:29]
  reg [34:0] sectored_entries_6_data_1; // @[TLB.scala 162:29]
  reg [34:0] sectored_entries_6_data_2; // @[TLB.scala 162:29]
  reg [34:0] sectored_entries_6_data_3; // @[TLB.scala 162:29]
  reg  sectored_entries_6_valid_0; // @[TLB.scala 162:29]
  reg  sectored_entries_6_valid_1; // @[TLB.scala 162:29]
  reg  sectored_entries_6_valid_2; // @[TLB.scala 162:29]
  reg  sectored_entries_6_valid_3; // @[TLB.scala 162:29]
  reg [26:0] sectored_entries_7_tag; // @[TLB.scala 162:29]
  reg [34:0] sectored_entries_7_data_0; // @[TLB.scala 162:29]
  reg [34:0] sectored_entries_7_data_1; // @[TLB.scala 162:29]
  reg [34:0] sectored_entries_7_data_2; // @[TLB.scala 162:29]
  reg [34:0] sectored_entries_7_data_3; // @[TLB.scala 162:29]
  reg  sectored_entries_7_valid_0; // @[TLB.scala 162:29]
  reg  sectored_entries_7_valid_1; // @[TLB.scala 162:29]
  reg  sectored_entries_7_valid_2; // @[TLB.scala 162:29]
  reg  sectored_entries_7_valid_3; // @[TLB.scala 162:29]
  reg [1:0] superpage_entries_0_level; // @[TLB.scala 163:30]
  reg [26:0] superpage_entries_0_tag; // @[TLB.scala 163:30]
  reg [34:0] superpage_entries_0_data_0; // @[TLB.scala 163:30]
  reg  superpage_entries_0_valid_0; // @[TLB.scala 163:30]
  reg [1:0] superpage_entries_1_level; // @[TLB.scala 163:30]
  reg [26:0] superpage_entries_1_tag; // @[TLB.scala 163:30]
  reg [34:0] superpage_entries_1_data_0; // @[TLB.scala 163:30]
  reg  superpage_entries_1_valid_0; // @[TLB.scala 163:30]
  reg [1:0] superpage_entries_2_level; // @[TLB.scala 163:30]
  reg [26:0] superpage_entries_2_tag; // @[TLB.scala 163:30]
  reg [34:0] superpage_entries_2_data_0; // @[TLB.scala 163:30]
  reg  superpage_entries_2_valid_0; // @[TLB.scala 163:30]
  reg [1:0] superpage_entries_3_level; // @[TLB.scala 163:30]
  reg [26:0] superpage_entries_3_tag; // @[TLB.scala 163:30]
  reg [34:0] superpage_entries_3_data_0; // @[TLB.scala 163:30]
  reg  superpage_entries_3_valid_0; // @[TLB.scala 163:30]
  reg [1:0] special_entry_level; // @[TLB.scala 164:56]
  reg [26:0] special_entry_tag; // @[TLB.scala 164:56]
  reg [34:0] special_entry_data_0; // @[TLB.scala 164:56]
  reg  special_entry_valid_0; // @[TLB.scala 164:56]
  reg [1:0] state; // @[TLB.scala 169:18]
  reg [26:0] r_refill_tag; // @[TLB.scala 170:25]
  reg [1:0] r_superpage_repl_addr; // @[TLB.scala 171:34]
  reg [2:0] r_sectored_repl_addr; // @[TLB.scala 172:33]
  reg [2:0] r_sectored_hit_addr; // @[TLB.scala 173:32]
  reg  r_sectored_hit; // @[TLB.scala 174:27]
  wire  priv_s = io_ptw_status_prv[0]; // @[TLB.scala 177:20]
  wire  priv_uses_vm = io_ptw_status_prv <= 2'h1; // @[TLB.scala 178:27]
  wire  vm_enabled = (io_ptw_ptbr_mode[3]) & priv_uses_vm; // @[TLB.scala 179:83]
  wire [26:0] vpn = io_req_bits_vaddr[38:12]; // @[TLB.scala 182:30]
  wire [19:0] refill_ppn = io_ptw_resp_bits_pte_ppn[19:0]; // @[TLB.scala 183:44]
  wire  _invalidate_refill_T = state == 2'h1; // @[package.scala 15:47]
  wire  _invalidate_refill_T_1 = state == 2'h3; // @[package.scala 15:47]
  wire  _invalidate_refill_T_2 = _invalidate_refill_T | _invalidate_refill_T_1; // @[package.scala 64:59]
  wire  invalidate_refill = _invalidate_refill_T_2 | io_sfence_valid; // @[TLB.scala 185:88]
  wire [1:0] mpu_ppn_right = mpu_ppn_data_barrier_io_y_ppn[19:18]; // @[TLB.scala 106:26]
  wire  mpu_ppn_ignore = special_entry_level < 2'h1; // @[TLB.scala 108:28]
  wire [26:0] _mpu_ppn_T_1 = mpu_ppn_ignore ? vpn : 27'h0; // @[TLB.scala 109:28]
  wire [26:0] _GEN_983 = {{7'd0}, mpu_ppn_data_barrier_io_y_ppn}; // @[TLB.scala 109:47]
  wire [26:0] _mpu_ppn_T_2 = _mpu_ppn_T_1 | _GEN_983; // @[TLB.scala 109:47]
  wire [8:0] mpu_ppn_left = _mpu_ppn_T_2[17:9]; // @[TLB.scala 109:58]
  wire  mpu_ppn_ignore_1 = special_entry_level < 2'h2; // @[TLB.scala 108:28]
  wire [26:0] _mpu_ppn_T_3 = mpu_ppn_ignore_1 ? vpn : 27'h0; // @[TLB.scala 109:28]
  wire [26:0] _mpu_ppn_T_4 = _mpu_ppn_T_3 | _GEN_983; // @[TLB.scala 109:47]
  wire [8:0] mpu_ppn_left_1 = _mpu_ppn_T_4[8:0]; // @[TLB.scala 109:58]
  wire [19:0] _mpu_ppn_T_5 = {mpu_ppn_right,mpu_ppn_left,mpu_ppn_left_1}; // @[Cat.scala 29:58]
  wire [27:0] _mpu_ppn_T_7 = vm_enabled ? {{8'd0}, _mpu_ppn_T_5} : io_req_bits_vaddr[39:12]; // @[TLB.scala 187:20]
  wire [27:0] mpu_ppn = io_ptw_resp_valid ? {{8'd0}, refill_ppn} : _mpu_ppn_T_7; // @[TLB.scala 186:20]
  wire [11:0] mpu_physaddr_left = io_req_bits_vaddr[11:0]; // @[TLB.scala 188:52]
  wire [39:0] mpu_physaddr = {mpu_ppn,mpu_physaddr_left}; // @[Cat.scala 29:58]
  wire [2:0] _mpu_priv_T_2 = {io_ptw_status_debug,io_ptw_status_prv}; // @[Cat.scala 29:58]
  wire [2:0] mpu_priv = io_ptw_resp_valid ? 3'h1 : _mpu_priv_T_2; // @[TLB.scala 189:27]
  wire [39:0] _legal_address_T = mpu_physaddr ^ 40'h3000; // @[Parameters.scala 138:31]
  wire [40:0] _legal_address_T_1 = {1'b0,$signed(_legal_address_T)}; // @[Parameters.scala 138:49]
  wire [40:0] _legal_address_T_3 = $signed(_legal_address_T_1) & -41'sh1000; // @[Parameters.scala 138:52]
  wire  _legal_address_T_4 = $signed(_legal_address_T_3) == 41'sh0; // @[Parameters.scala 138:67]
  wire [39:0] _legal_address_T_5 = mpu_physaddr ^ 40'hc000000; // @[Parameters.scala 138:31]
  wire [40:0] _legal_address_T_6 = {1'b0,$signed(_legal_address_T_5)}; // @[Parameters.scala 138:49]
  wire [40:0] _legal_address_T_8 = $signed(_legal_address_T_6) & -41'sh4000000; // @[Parameters.scala 138:52]
  wire  _legal_address_T_9 = $signed(_legal_address_T_8) == 41'sh0; // @[Parameters.scala 138:67]
  wire [39:0] _legal_address_T_10 = mpu_physaddr ^ 40'h2000000; // @[Parameters.scala 138:31]
  wire [40:0] _legal_address_T_11 = {1'b0,$signed(_legal_address_T_10)}; // @[Parameters.scala 138:49]
  wire [40:0] _legal_address_T_13 = $signed(_legal_address_T_11) & -41'sh10000; // @[Parameters.scala 138:52]
  wire  _legal_address_T_14 = $signed(_legal_address_T_13) == 41'sh0; // @[Parameters.scala 138:67]
  wire [40:0] _legal_address_T_16 = {1'b0,$signed(mpu_physaddr)}; // @[Parameters.scala 138:49]
  wire [40:0] _legal_address_T_18 = $signed(_legal_address_T_16) & -41'sh1000; // @[Parameters.scala 138:52]
  wire  _legal_address_T_19 = $signed(_legal_address_T_18) == 41'sh0; // @[Parameters.scala 138:67]
  wire [39:0] _legal_address_T_20 = mpu_physaddr ^ 40'h10000; // @[Parameters.scala 138:31]
  wire [40:0] _legal_address_T_21 = {1'b0,$signed(_legal_address_T_20)}; // @[Parameters.scala 138:49]
  wire [40:0] _legal_address_T_23 = $signed(_legal_address_T_21) & -41'sh10000; // @[Parameters.scala 138:52]
  wire  _legal_address_T_24 = $signed(_legal_address_T_23) == 41'sh0; // @[Parameters.scala 138:67]
  wire [39:0] _legal_address_T_25 = mpu_physaddr ^ 40'h80000000; // @[Parameters.scala 138:31]
  wire [40:0] _legal_address_T_26 = {1'b0,$signed(_legal_address_T_25)}; // @[Parameters.scala 138:49]
  wire [40:0] _legal_address_T_28 = $signed(_legal_address_T_26) & -41'sh10000000; // @[Parameters.scala 138:52]
  wire  _legal_address_T_29 = $signed(_legal_address_T_28) == 41'sh0; // @[Parameters.scala 138:67]
  wire [39:0] _legal_address_T_30 = mpu_physaddr ^ 40'h60000000; // @[Parameters.scala 138:31]
  wire [40:0] _legal_address_T_31 = {1'b0,$signed(_legal_address_T_30)}; // @[Parameters.scala 138:49]
  wire [40:0] _legal_address_T_33 = $signed(_legal_address_T_31) & -41'sh20000000; // @[Parameters.scala 138:52]
  wire  _legal_address_T_34 = $signed(_legal_address_T_33) == 41'sh0; // @[Parameters.scala 138:67]
  wire  legal_address = (((((_legal_address_T_4 | _legal_address_T_9) | _legal_address_T_14) | _legal_address_T_19) |
    _legal_address_T_24) | _legal_address_T_29) | _legal_address_T_34; // @[TLB.scala 195:67]
  wire [40:0] _cacheable_T_8 = $signed(_legal_address_T_26) & 41'sh80000000; // @[Parameters.scala 138:52]
  wire  _cacheable_T_9 = $signed(_cacheable_T_8) == 41'sh0; // @[Parameters.scala 138:67]
  wire  cacheable = legal_address & _cacheable_T_9; // @[TLB.scala 197:19]
  wire [39:0] _homogeneous_T_54 = mpu_physaddr ^ 40'h8000000; // @[Parameters.scala 138:31]
  wire [40:0] _homogeneous_T_55 = {1'b0,$signed(_homogeneous_T_54)}; // @[Parameters.scala 138:49]
  wire [40:0] _homogeneous_T_57 = $signed(_homogeneous_T_55) & 41'shc8000000; // @[Parameters.scala 138:52]
  wire  _homogeneous_T_58 = $signed(_homogeneous_T_57) == 41'sh0; // @[Parameters.scala 138:67]
  wire [40:0] _homogeneous_T_71 = $signed(_legal_address_T_16) & 41'shc8010000; // @[Parameters.scala 138:52]
  wire  _homogeneous_T_72 = $signed(_homogeneous_T_71) == 41'sh0; // @[Parameters.scala 138:67]
  wire  _homogeneous_T_79 = _homogeneous_T_72 | _homogeneous_T_58; // @[TLBPermissions.scala 82:66]
  wire  deny_access_to_debug = (mpu_priv <= 3'h3) & _legal_address_T_19; // @[TLB.scala 200:48]
  wire  _prot_r_T_6 = ~deny_access_to_debug; // @[TLB.scala 201:44]
  wire  prot_r = (legal_address & (~deny_access_to_debug)) & pmp_io_r; // @[TLB.scala 201:66]
  wire [39:0] _prot_w_T_10 = mpu_physaddr ^ 40'h40000000; // @[Parameters.scala 138:31]
  wire [40:0] _prot_w_T_11 = {1'b0,$signed(_prot_w_T_10)}; // @[Parameters.scala 138:49]
  wire [40:0] _prot_w_T_13 = $signed(_prot_w_T_11) & 41'shc0000000; // @[Parameters.scala 138:52]
  wire  _prot_w_T_14 = $signed(_prot_w_T_13) == 41'sh0; // @[Parameters.scala 138:67]
  wire [40:0] _prot_w_T_18 = $signed(_legal_address_T_26) & 41'shc0000000; // @[Parameters.scala 138:52]
  wire  _prot_w_T_19 = $signed(_prot_w_T_18) == 41'sh0; // @[Parameters.scala 138:67]
  wire  _prot_w_T_22 = (_homogeneous_T_79 | _prot_w_T_14) | _prot_w_T_19; // @[Parameters.scala 616:89]
  wire  _prot_w_T_31 = legal_address & _prot_w_T_22; // @[TLB.scala 197:19]
  wire  prot_w = (_prot_w_T_31 & _prot_r_T_6) & pmp_io_w; // @[TLB.scala 202:70]
  wire  prot_al = legal_address & _homogeneous_T_79; // @[TLB.scala 197:19]
  wire [40:0] _prot_x_T_3 = $signed(_legal_address_T_16) & 41'shca000000; // @[Parameters.scala 138:52]
  wire  _prot_x_T_4 = $signed(_prot_x_T_3) == 41'sh0; // @[Parameters.scala 138:67]
  wire  _prot_x_T_16 = (_prot_x_T_4 | _prot_w_T_14) | _prot_w_T_19; // @[Parameters.scala 616:89]
  wire  _prot_x_T_31 = legal_address & _prot_x_T_16; // @[TLB.scala 197:19]
  wire  prot_x = (_prot_x_T_31 & _prot_r_T_6) & pmp_io_x; // @[TLB.scala 206:65]
  wire [40:0] _prot_eff_T_20 = $signed(_legal_address_T_16) & 41'shca012000; // @[Parameters.scala 138:52]
  wire  _prot_eff_T_21 = $signed(_prot_eff_T_20) == 41'sh0; // @[Parameters.scala 138:67]
  wire [40:0] _prot_eff_T_25 = $signed(_legal_address_T_11) & 41'shca010000; // @[Parameters.scala 138:52]
  wire  _prot_eff_T_26 = $signed(_prot_eff_T_25) == 41'sh0; // @[Parameters.scala 138:67]
  wire  _prot_eff_T_39 = ((_prot_eff_T_21 | _prot_eff_T_26) | _homogeneous_T_58) | _prot_w_T_14; // @[Parameters.scala 616:89]
  wire  prot_eff = legal_address & _prot_eff_T_39; // @[TLB.scala 197:19]
  wire  _sector_hits_T_2 = ((sectored_entries_0_valid_0 | sectored_entries_0_valid_1) | sectored_entries_0_valid_2) |
    sectored_entries_0_valid_3; // @[package.scala 64:59]
  wire [26:0] _sector_hits_T_3 = sectored_entries_0_tag ^ vpn; // @[TLB.scala 88:41]
  wire  _sector_hits_T_5 = (_sector_hits_T_3[26:2]) == 25'h0; // @[TLB.scala 88:66]
  wire  sector_hits_0 = _sector_hits_T_2 & _sector_hits_T_5; // @[TLB.scala 87:40]
  wire  _sector_hits_T_8 = ((sectored_entries_1_valid_0 | sectored_entries_1_valid_1) | sectored_entries_1_valid_2) |
    sectored_entries_1_valid_3; // @[package.scala 64:59]
  wire [26:0] _sector_hits_T_9 = sectored_entries_1_tag ^ vpn; // @[TLB.scala 88:41]
  wire  _sector_hits_T_11 = (_sector_hits_T_9[26:2]) == 25'h0; // @[TLB.scala 88:66]
  wire  sector_hits_1 = _sector_hits_T_8 & _sector_hits_T_11; // @[TLB.scala 87:40]
  wire  _sector_hits_T_14 = ((sectored_entries_2_valid_0 | sectored_entries_2_valid_1) | sectored_entries_2_valid_2) |
    sectored_entries_2_valid_3; // @[package.scala 64:59]
  wire [26:0] _sector_hits_T_15 = sectored_entries_2_tag ^ vpn; // @[TLB.scala 88:41]
  wire  _sector_hits_T_17 = (_sector_hits_T_15[26:2]) == 25'h0; // @[TLB.scala 88:66]
  wire  sector_hits_2 = _sector_hits_T_14 & _sector_hits_T_17; // @[TLB.scala 87:40]
  wire  _sector_hits_T_20 = ((sectored_entries_3_valid_0 | sectored_entries_3_valid_1) | sectored_entries_3_valid_2) |
    sectored_entries_3_valid_3; // @[package.scala 64:59]
  wire [26:0] _sector_hits_T_21 = sectored_entries_3_tag ^ vpn; // @[TLB.scala 88:41]
  wire  _sector_hits_T_23 = (_sector_hits_T_21[26:2]) == 25'h0; // @[TLB.scala 88:66]
  wire  sector_hits_3 = _sector_hits_T_20 & _sector_hits_T_23; // @[TLB.scala 87:40]
  wire  _sector_hits_T_26 = ((sectored_entries_4_valid_0 | sectored_entries_4_valid_1) | sectored_entries_4_valid_2) |
    sectored_entries_4_valid_3; // @[package.scala 64:59]
  wire [26:0] _sector_hits_T_27 = sectored_entries_4_tag ^ vpn; // @[TLB.scala 88:41]
  wire  _sector_hits_T_29 = (_sector_hits_T_27[26:2]) == 25'h0; // @[TLB.scala 88:66]
  wire  sector_hits_4 = _sector_hits_T_26 & _sector_hits_T_29; // @[TLB.scala 87:40]
  wire  _sector_hits_T_32 = ((sectored_entries_5_valid_0 | sectored_entries_5_valid_1) | sectored_entries_5_valid_2) |
    sectored_entries_5_valid_3; // @[package.scala 64:59]
  wire [26:0] _sector_hits_T_33 = sectored_entries_5_tag ^ vpn; // @[TLB.scala 88:41]
  wire  _sector_hits_T_35 = (_sector_hits_T_33[26:2]) == 25'h0; // @[TLB.scala 88:66]
  wire  sector_hits_5 = _sector_hits_T_32 & _sector_hits_T_35; // @[TLB.scala 87:40]
  wire  _sector_hits_T_38 = ((sectored_entries_6_valid_0 | sectored_entries_6_valid_1) | sectored_entries_6_valid_2) |
    sectored_entries_6_valid_3; // @[package.scala 64:59]
  wire [26:0] _sector_hits_T_39 = sectored_entries_6_tag ^ vpn; // @[TLB.scala 88:41]
  wire  _sector_hits_T_41 = (_sector_hits_T_39[26:2]) == 25'h0; // @[TLB.scala 88:66]
  wire  sector_hits_6 = _sector_hits_T_38 & _sector_hits_T_41; // @[TLB.scala 87:40]
  wire  _sector_hits_T_44 = ((sectored_entries_7_valid_0 | sectored_entries_7_valid_1) | sectored_entries_7_valid_2) |
    sectored_entries_7_valid_3; // @[package.scala 64:59]
  wire [26:0] _sector_hits_T_45 = sectored_entries_7_tag ^ vpn; // @[TLB.scala 88:41]
  wire  _sector_hits_T_47 = (_sector_hits_T_45[26:2]) == 25'h0; // @[TLB.scala 88:66]
  wire  sector_hits_7 = _sector_hits_T_44 & _sector_hits_T_47; // @[TLB.scala 87:40]
  wire  superpage_hits_ignore_1 = superpage_entries_0_level < 2'h1; // @[TLB.scala 94:28]
  wire  superpage_hits_0 = (superpage_entries_0_valid_0 & ((superpage_entries_0_tag[26:18]) == (vpn[26:18]))) & (
    superpage_hits_ignore_1 | ((superpage_entries_0_tag[17:9]) == (vpn[17:9]))); // @[TLB.scala 95:29]
  wire  superpage_hits_ignore_4 = superpage_entries_1_level < 2'h1; // @[TLB.scala 94:28]
  wire  superpage_hits_1 = (superpage_entries_1_valid_0 & ((superpage_entries_1_tag[26:18]) == (vpn[26:18]))) & (
    superpage_hits_ignore_4 | ((superpage_entries_1_tag[17:9]) == (vpn[17:9]))); // @[TLB.scala 95:29]
  wire  superpage_hits_ignore_7 = superpage_entries_2_level < 2'h1; // @[TLB.scala 94:28]
  wire  superpage_hits_2 = (superpage_entries_2_valid_0 & ((superpage_entries_2_tag[26:18]) == (vpn[26:18]))) & (
    superpage_hits_ignore_7 | ((superpage_entries_2_tag[17:9]) == (vpn[17:9]))); // @[TLB.scala 95:29]
  wire  superpage_hits_ignore_10 = superpage_entries_3_level < 2'h1; // @[TLB.scala 94:28]
  wire  superpage_hits_3 = (superpage_entries_3_valid_0 & ((superpage_entries_3_tag[26:18]) == (vpn[26:18]))) & (
    superpage_hits_ignore_10 | ((superpage_entries_3_tag[17:9]) == (vpn[17:9]))); // @[TLB.scala 95:29]
  wire [1:0] hitsVec_idx = vpn[1:0]; // @[package.scala 143:13]
  wire  _GEN_1 = 2'h1 == hitsVec_idx ? sectored_entries_0_valid_1 : sectored_entries_0_valid_0; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  _GEN_2 = 2'h2 == hitsVec_idx ? sectored_entries_0_valid_2 : _GEN_1; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  _GEN_3 = 2'h3 == hitsVec_idx ? sectored_entries_0_valid_3 : _GEN_2; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  _hitsVec_T_3 = _GEN_3 & _sector_hits_T_5; // @[TLB.scala 100:18]
  wire  hitsVec_0 = vm_enabled & _hitsVec_T_3; // @[TLB.scala 211:44]
  wire  _GEN_5 = 2'h1 == hitsVec_idx ? sectored_entries_1_valid_1 : sectored_entries_1_valid_0; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  _GEN_6 = 2'h2 == hitsVec_idx ? sectored_entries_1_valid_2 : _GEN_5; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  _GEN_7 = 2'h3 == hitsVec_idx ? sectored_entries_1_valid_3 : _GEN_6; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  _hitsVec_T_7 = _GEN_7 & _sector_hits_T_11; // @[TLB.scala 100:18]
  wire  hitsVec_1 = vm_enabled & _hitsVec_T_7; // @[TLB.scala 211:44]
  wire  _GEN_9 = 2'h1 == hitsVec_idx ? sectored_entries_2_valid_1 : sectored_entries_2_valid_0; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  _GEN_10 = 2'h2 == hitsVec_idx ? sectored_entries_2_valid_2 : _GEN_9; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  _GEN_11 = 2'h3 == hitsVec_idx ? sectored_entries_2_valid_3 : _GEN_10; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  _hitsVec_T_11 = _GEN_11 & _sector_hits_T_17; // @[TLB.scala 100:18]
  wire  hitsVec_2 = vm_enabled & _hitsVec_T_11; // @[TLB.scala 211:44]
  wire  _GEN_13 = 2'h1 == hitsVec_idx ? sectored_entries_3_valid_1 : sectored_entries_3_valid_0; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  _GEN_14 = 2'h2 == hitsVec_idx ? sectored_entries_3_valid_2 : _GEN_13; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  _GEN_15 = 2'h3 == hitsVec_idx ? sectored_entries_3_valid_3 : _GEN_14; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  _hitsVec_T_15 = _GEN_15 & _sector_hits_T_23; // @[TLB.scala 100:18]
  wire  hitsVec_3 = vm_enabled & _hitsVec_T_15; // @[TLB.scala 211:44]
  wire  _GEN_17 = 2'h1 == hitsVec_idx ? sectored_entries_4_valid_1 : sectored_entries_4_valid_0; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  _GEN_18 = 2'h2 == hitsVec_idx ? sectored_entries_4_valid_2 : _GEN_17; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  _GEN_19 = 2'h3 == hitsVec_idx ? sectored_entries_4_valid_3 : _GEN_18; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  _hitsVec_T_19 = _GEN_19 & _sector_hits_T_29; // @[TLB.scala 100:18]
  wire  hitsVec_4 = vm_enabled & _hitsVec_T_19; // @[TLB.scala 211:44]
  wire  _GEN_21 = 2'h1 == hitsVec_idx ? sectored_entries_5_valid_1 : sectored_entries_5_valid_0; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  _GEN_22 = 2'h2 == hitsVec_idx ? sectored_entries_5_valid_2 : _GEN_21; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  _GEN_23 = 2'h3 == hitsVec_idx ? sectored_entries_5_valid_3 : _GEN_22; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  _hitsVec_T_23 = _GEN_23 & _sector_hits_T_35; // @[TLB.scala 100:18]
  wire  hitsVec_5 = vm_enabled & _hitsVec_T_23; // @[TLB.scala 211:44]
  wire  _GEN_25 = 2'h1 == hitsVec_idx ? sectored_entries_6_valid_1 : sectored_entries_6_valid_0; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  _GEN_26 = 2'h2 == hitsVec_idx ? sectored_entries_6_valid_2 : _GEN_25; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  _GEN_27 = 2'h3 == hitsVec_idx ? sectored_entries_6_valid_3 : _GEN_26; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  _hitsVec_T_27 = _GEN_27 & _sector_hits_T_41; // @[TLB.scala 100:18]
  wire  hitsVec_6 = vm_enabled & _hitsVec_T_27; // @[TLB.scala 211:44]
  wire  _GEN_29 = 2'h1 == hitsVec_idx ? sectored_entries_7_valid_1 : sectored_entries_7_valid_0; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  _GEN_30 = 2'h2 == hitsVec_idx ? sectored_entries_7_valid_2 : _GEN_29; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  _GEN_31 = 2'h3 == hitsVec_idx ? sectored_entries_7_valid_3 : _GEN_30; // @[TLB.scala 100:18 TLB.scala 100:18]
  wire  _hitsVec_T_31 = _GEN_31 & _sector_hits_T_47; // @[TLB.scala 100:18]
  wire  hitsVec_7 = vm_enabled & _hitsVec_T_31; // @[TLB.scala 211:44]
  wire  hitsVec_8 = vm_enabled & superpage_hits_0; // @[TLB.scala 211:44]
  wire  hitsVec_9 = vm_enabled & superpage_hits_1; // @[TLB.scala 211:44]
  wire  hitsVec_10 = vm_enabled & superpage_hits_2; // @[TLB.scala 211:44]
  wire  hitsVec_11 = vm_enabled & superpage_hits_3; // @[TLB.scala 211:44]
  wire  _hitsVec_T_106 = ((special_entry_valid_0 & ((special_entry_tag[26:18]) == (vpn[26:18]))) & (mpu_ppn_ignore | ((
    special_entry_tag[17:9]) == (vpn[17:9])))) & (mpu_ppn_ignore_1 | ((special_entry_tag[8:0]) == (vpn[8:0]))); // @[TLB.scala 95:29]
  wire  hitsVec_12 = vm_enabled & _hitsVec_T_106; // @[TLB.scala 211:44]
  wire [5:0] real_hits_left = {hitsVec_5,hitsVec_4,hitsVec_3,hitsVec_2,hitsVec_1,hitsVec_0}; // @[Cat.scala 29:58]
  wire [12:0] real_hits = {hitsVec_12,hitsVec_11,hitsVec_10,hitsVec_9,hitsVec_8,hitsVec_7,hitsVec_6,real_hits_left}; // @[Cat.scala 29:58]
  wire  hits_right = ~vm_enabled; // @[TLB.scala 213:18]
  wire [13:0] hits = {hits_right,hitsVec_12,hitsVec_11,hitsVec_10,hitsVec_9,hitsVec_8,hitsVec_7,hitsVec_6,real_hits_left
    }; // @[Cat.scala 29:58]
  wire [34:0] _GEN_33 = 2'h1 == hitsVec_idx ? sectored_entries_0_data_1 : sectored_entries_0_data_0; // @[]
  wire [34:0] _GEN_34 = 2'h2 == hitsVec_idx ? sectored_entries_0_data_2 : _GEN_33; // @[]
  wire [34:0] _GEN_35 = 2'h3 == hitsVec_idx ? sectored_entries_0_data_3 : _GEN_34; // @[]
  wire [34:0] _GEN_37 = 2'h1 == hitsVec_idx ? sectored_entries_1_data_1 : sectored_entries_1_data_0; // @[]
  wire [34:0] _GEN_38 = 2'h2 == hitsVec_idx ? sectored_entries_1_data_2 : _GEN_37; // @[]
  wire [34:0] _GEN_39 = 2'h3 == hitsVec_idx ? sectored_entries_1_data_3 : _GEN_38; // @[]
  wire [34:0] _GEN_41 = 2'h1 == hitsVec_idx ? sectored_entries_2_data_1 : sectored_entries_2_data_0; // @[]
  wire [34:0] _GEN_42 = 2'h2 == hitsVec_idx ? sectored_entries_2_data_2 : _GEN_41; // @[]
  wire [34:0] _GEN_43 = 2'h3 == hitsVec_idx ? sectored_entries_2_data_3 : _GEN_42; // @[]
  wire [34:0] _GEN_45 = 2'h1 == hitsVec_idx ? sectored_entries_3_data_1 : sectored_entries_3_data_0; // @[]
  wire [34:0] _GEN_46 = 2'h2 == hitsVec_idx ? sectored_entries_3_data_2 : _GEN_45; // @[]
  wire [34:0] _GEN_47 = 2'h3 == hitsVec_idx ? sectored_entries_3_data_3 : _GEN_46; // @[]
  wire [34:0] _GEN_49 = 2'h1 == hitsVec_idx ? sectored_entries_4_data_1 : sectored_entries_4_data_0; // @[]
  wire [34:0] _GEN_50 = 2'h2 == hitsVec_idx ? sectored_entries_4_data_2 : _GEN_49; // @[]
  wire [34:0] _GEN_51 = 2'h3 == hitsVec_idx ? sectored_entries_4_data_3 : _GEN_50; // @[]
  wire [34:0] _GEN_53 = 2'h1 == hitsVec_idx ? sectored_entries_5_data_1 : sectored_entries_5_data_0; // @[]
  wire [34:0] _GEN_54 = 2'h2 == hitsVec_idx ? sectored_entries_5_data_2 : _GEN_53; // @[]
  wire [34:0] _GEN_55 = 2'h3 == hitsVec_idx ? sectored_entries_5_data_3 : _GEN_54; // @[]
  wire [34:0] _GEN_57 = 2'h1 == hitsVec_idx ? sectored_entries_6_data_1 : sectored_entries_6_data_0; // @[]
  wire [34:0] _GEN_58 = 2'h2 == hitsVec_idx ? sectored_entries_6_data_2 : _GEN_57; // @[]
  wire [34:0] _GEN_59 = 2'h3 == hitsVec_idx ? sectored_entries_6_data_3 : _GEN_58; // @[]
  wire [34:0] _GEN_61 = 2'h1 == hitsVec_idx ? sectored_entries_7_data_1 : sectored_entries_7_data_0; // @[]
  wire [34:0] _GEN_62 = 2'h2 == hitsVec_idx ? sectored_entries_7_data_2 : _GEN_61; // @[]
  wire [34:0] _GEN_63 = 2'h3 == hitsVec_idx ? sectored_entries_7_data_3 : _GEN_62; // @[]
  wire [1:0] ppn_right = ppn_data_barrier_8_io_y_ppn[19:18]; // @[TLB.scala 106:26]
  wire [26:0] _ppn_T_1 = superpage_hits_ignore_1 ? vpn : 27'h0; // @[TLB.scala 109:28]
  wire [26:0] _GEN_985 = {{7'd0}, ppn_data_barrier_8_io_y_ppn}; // @[TLB.scala 109:47]
  wire [26:0] _ppn_T_2 = _ppn_T_1 | _GEN_985; // @[TLB.scala 109:47]
  wire [8:0] ppn_left = _ppn_T_2[17:9]; // @[TLB.scala 109:58]
  wire [26:0] _ppn_T_4 = vpn | _GEN_985; // @[TLB.scala 109:47]
  wire [8:0] ppn_left_1 = _ppn_T_4[8:0]; // @[TLB.scala 109:58]
  wire [19:0] _ppn_T_5 = {ppn_right,ppn_left,ppn_left_1}; // @[Cat.scala 29:58]
  wire [1:0] ppn_right_2 = ppn_data_barrier_9_io_y_ppn[19:18]; // @[TLB.scala 106:26]
  wire [26:0] _ppn_T_6 = superpage_hits_ignore_4 ? vpn : 27'h0; // @[TLB.scala 109:28]
  wire [26:0] _GEN_987 = {{7'd0}, ppn_data_barrier_9_io_y_ppn}; // @[TLB.scala 109:47]
  wire [26:0] _ppn_T_7 = _ppn_T_6 | _GEN_987; // @[TLB.scala 109:47]
  wire [8:0] ppn_left_2 = _ppn_T_7[17:9]; // @[TLB.scala 109:58]
  wire [26:0] _ppn_T_9 = vpn | _GEN_987; // @[TLB.scala 109:47]
  wire [8:0] ppn_left_3 = _ppn_T_9[8:0]; // @[TLB.scala 109:58]
  wire [19:0] _ppn_T_10 = {ppn_right_2,ppn_left_2,ppn_left_3}; // @[Cat.scala 29:58]
  wire [1:0] ppn_right_4 = ppn_data_barrier_10_io_y_ppn[19:18]; // @[TLB.scala 106:26]
  wire [26:0] _ppn_T_11 = superpage_hits_ignore_7 ? vpn : 27'h0; // @[TLB.scala 109:28]
  wire [26:0] _GEN_989 = {{7'd0}, ppn_data_barrier_10_io_y_ppn}; // @[TLB.scala 109:47]
  wire [26:0] _ppn_T_12 = _ppn_T_11 | _GEN_989; // @[TLB.scala 109:47]
  wire [8:0] ppn_left_4 = _ppn_T_12[17:9]; // @[TLB.scala 109:58]
  wire [26:0] _ppn_T_14 = vpn | _GEN_989; // @[TLB.scala 109:47]
  wire [8:0] ppn_left_5 = _ppn_T_14[8:0]; // @[TLB.scala 109:58]
  wire [19:0] _ppn_T_15 = {ppn_right_4,ppn_left_4,ppn_left_5}; // @[Cat.scala 29:58]
  wire [1:0] ppn_right_6 = ppn_data_barrier_11_io_y_ppn[19:18]; // @[TLB.scala 106:26]
  wire [26:0] _ppn_T_16 = superpage_hits_ignore_10 ? vpn : 27'h0; // @[TLB.scala 109:28]
  wire [26:0] _GEN_991 = {{7'd0}, ppn_data_barrier_11_io_y_ppn}; // @[TLB.scala 109:47]
  wire [26:0] _ppn_T_17 = _ppn_T_16 | _GEN_991; // @[TLB.scala 109:47]
  wire [8:0] ppn_left_6 = _ppn_T_17[17:9]; // @[TLB.scala 109:58]
  wire [26:0] _ppn_T_19 = vpn | _GEN_991; // @[TLB.scala 109:47]
  wire [8:0] ppn_left_7 = _ppn_T_19[8:0]; // @[TLB.scala 109:58]
  wire [19:0] _ppn_T_20 = {ppn_right_6,ppn_left_6,ppn_left_7}; // @[Cat.scala 29:58]
  wire [1:0] ppn_right_8 = ppn_data_barrier_12_io_y_ppn[19:18]; // @[TLB.scala 106:26]
  wire [26:0] _GEN_993 = {{7'd0}, ppn_data_barrier_12_io_y_ppn}; // @[TLB.scala 109:47]
  wire [26:0] _ppn_T_22 = _mpu_ppn_T_1 | _GEN_993; // @[TLB.scala 109:47]
  wire [8:0] ppn_left_8 = _ppn_T_22[17:9]; // @[TLB.scala 109:58]
  wire [26:0] _ppn_T_24 = _mpu_ppn_T_3 | _GEN_993; // @[TLB.scala 109:47]
  wire [8:0] ppn_left_9 = _ppn_T_24[8:0]; // @[TLB.scala 109:58]
  wire [19:0] _ppn_T_25 = {ppn_right_8,ppn_left_8,ppn_left_9}; // @[Cat.scala 29:58]
  wire [19:0] _ppn_T_27 = hitsVec_0 ? ppn_data_barrier_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_28 = hitsVec_1 ? ppn_data_barrier_1_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_29 = hitsVec_2 ? ppn_data_barrier_2_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_30 = hitsVec_3 ? ppn_data_barrier_3_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_31 = hitsVec_4 ? ppn_data_barrier_4_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_32 = hitsVec_5 ? ppn_data_barrier_5_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_33 = hitsVec_6 ? ppn_data_barrier_6_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_34 = hitsVec_7 ? ppn_data_barrier_7_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_35 = hitsVec_8 ? _ppn_T_5 : 20'h0; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_36 = hitsVec_9 ? _ppn_T_10 : 20'h0; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_37 = hitsVec_10 ? _ppn_T_15 : 20'h0; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_38 = hitsVec_11 ? _ppn_T_20 : 20'h0; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_39 = hitsVec_12 ? _ppn_T_25 : 20'h0; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_40 = hits_right ? vpn[19:0] : 20'h0; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_41 = _ppn_T_27 | _ppn_T_28; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_42 = _ppn_T_41 | _ppn_T_29; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_43 = _ppn_T_42 | _ppn_T_30; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_44 = _ppn_T_43 | _ppn_T_31; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_45 = _ppn_T_44 | _ppn_T_32; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_46 = _ppn_T_45 | _ppn_T_33; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_47 = _ppn_T_46 | _ppn_T_34; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_48 = _ppn_T_47 | _ppn_T_35; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_49 = _ppn_T_48 | _ppn_T_36; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_50 = _ppn_T_49 | _ppn_T_37; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_51 = _ppn_T_50 | _ppn_T_38; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_52 = _ppn_T_51 | _ppn_T_39; // @[Mux.scala 27:72]
  wire [19:0] ppn = _ppn_T_52 | _ppn_T_40; // @[Mux.scala 27:72]
  wire  newEntry_g = io_ptw_resp_bits_pte_g & io_ptw_resp_bits_pte_v; // @[TLB.scala 223:25]
  wire  _newEntry_sr_T_4 = (io_ptw_resp_bits_pte_v & (io_ptw_resp_bits_pte_r | (io_ptw_resp_bits_pte_x & (~
    io_ptw_resp_bits_pte_w)))) & io_ptw_resp_bits_pte_a; // @[PTW.scala 70:52]
  wire  newEntry_sr = _newEntry_sr_T_4 & io_ptw_resp_bits_pte_r; // @[PTW.scala 74:35]
  wire  newEntry_sw = (_newEntry_sr_T_4 & io_ptw_resp_bits_pte_w) & io_ptw_resp_bits_pte_d; // @[PTW.scala 75:40]
  wire  newEntry_sx = _newEntry_sr_T_4 & io_ptw_resp_bits_pte_x; // @[PTW.scala 76:35]
  wire  _T = ~io_ptw_resp_bits_homogeneous; // @[TLB.scala 237:37]
  wire [7:0] special_entry_data_0_left = {prot_x,prot_r,_prot_w_T_31,prot_al,prot_al,prot_eff,cacheable,1'h0}; // @[TLB.scala 123:24]
  wire [34:0] _special_entry_data_0_T = {refill_ppn,io_ptw_resp_bits_pte_u,newEntry_g,io_ptw_resp_bits_ae,newEntry_sw,
    newEntry_sx,newEntry_sr,prot_w,special_entry_data_0_left}; // @[TLB.scala 123:24]
  wire  _GEN_64 = invalidate_refill ? 1'h0 : 1'h1; // @[TLB.scala 240:34 TLB.scala 126:38 TLB.scala 122:16]
  wire  _T_2 = io_ptw_resp_bits_level < 2'h2; // @[TLB.scala 242:40]
  wire  _T_3 = r_superpage_repl_addr == 2'h0; // @[TLB.scala 243:82]
  wire  _GEN_67 = _T_3 ? _GEN_64 : superpage_entries_0_valid_0; // @[TLB.scala 243:89 TLB.scala 163:30]
  wire  _T_4 = r_superpage_repl_addr == 2'h1; // @[TLB.scala 243:82]
  wire  _GEN_71 = _T_4 ? _GEN_64 : superpage_entries_1_valid_0; // @[TLB.scala 243:89 TLB.scala 163:30]
  wire  _T_5 = r_superpage_repl_addr == 2'h2; // @[TLB.scala 243:82]
  wire  _GEN_75 = _T_5 ? _GEN_64 : superpage_entries_2_valid_0; // @[TLB.scala 243:89 TLB.scala 163:30]
  wire  _T_6 = r_superpage_repl_addr == 2'h3; // @[TLB.scala 243:82]
  wire  _GEN_79 = _T_6 ? _GEN_64 : superpage_entries_3_valid_0; // @[TLB.scala 243:89 TLB.scala 163:30]
  wire [2:0] waddr = r_sectored_hit ? r_sectored_hit_addr : r_sectored_repl_addr; // @[TLB.scala 248:22]
  wire  _T_7 = waddr == 3'h0; // @[TLB.scala 249:65]
  wire  _T_8 = ~r_sectored_hit; // @[TLB.scala 250:15]
  wire  _GEN_81 = _T_8 ? 1'h0 : sectored_entries_0_valid_0; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  _GEN_82 = _T_8 ? 1'h0 : sectored_entries_0_valid_1; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  _GEN_83 = _T_8 ? 1'h0 : sectored_entries_0_valid_2; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  _GEN_84 = _T_8 ? 1'h0 : sectored_entries_0_valid_3; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire [1:0] idx = r_refill_tag[1:0]; // @[package.scala 143:13]
  wire  _GEN_85 = (2'h0 == idx) | _GEN_81; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  _GEN_86 = (2'h1 == idx) | _GEN_82; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  _GEN_87 = (2'h2 == idx) | _GEN_83; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  _GEN_88 = (2'h3 == idx) | _GEN_84; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire [34:0] _GEN_89 = 2'h0 == idx ? _special_entry_data_0_T : sectored_entries_0_data_0; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] _GEN_90 = 2'h1 == idx ? _special_entry_data_0_T : sectored_entries_0_data_1; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] _GEN_91 = 2'h2 == idx ? _special_entry_data_0_T : sectored_entries_0_data_2; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] _GEN_92 = 2'h3 == idx ? _special_entry_data_0_T : sectored_entries_0_data_3; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire  _GEN_93 = invalidate_refill ? 1'h0 : _GEN_85; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  _GEN_94 = invalidate_refill ? 1'h0 : _GEN_86; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  _GEN_95 = invalidate_refill ? 1'h0 : _GEN_87; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  _GEN_96 = invalidate_refill ? 1'h0 : _GEN_88; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  _GEN_97 = _T_7 ? _GEN_93 : sectored_entries_0_valid_0; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  _GEN_98 = _T_7 ? _GEN_94 : sectored_entries_0_valid_1; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  _GEN_99 = _T_7 ? _GEN_95 : sectored_entries_0_valid_2; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  _GEN_100 = _T_7 ? _GEN_96 : sectored_entries_0_valid_3; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  _T_9 = waddr == 3'h1; // @[TLB.scala 249:65]
  wire  _GEN_107 = _T_8 ? 1'h0 : sectored_entries_1_valid_0; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  _GEN_108 = _T_8 ? 1'h0 : sectored_entries_1_valid_1; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  _GEN_109 = _T_8 ? 1'h0 : sectored_entries_1_valid_2; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  _GEN_110 = _T_8 ? 1'h0 : sectored_entries_1_valid_3; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  _GEN_111 = (2'h0 == idx) | _GEN_107; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  _GEN_112 = (2'h1 == idx) | _GEN_108; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  _GEN_113 = (2'h2 == idx) | _GEN_109; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  _GEN_114 = (2'h3 == idx) | _GEN_110; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire [34:0] _GEN_115 = 2'h0 == idx ? _special_entry_data_0_T : sectored_entries_1_data_0; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] _GEN_116 = 2'h1 == idx ? _special_entry_data_0_T : sectored_entries_1_data_1; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] _GEN_117 = 2'h2 == idx ? _special_entry_data_0_T : sectored_entries_1_data_2; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] _GEN_118 = 2'h3 == idx ? _special_entry_data_0_T : sectored_entries_1_data_3; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire  _GEN_119 = invalidate_refill ? 1'h0 : _GEN_111; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  _GEN_120 = invalidate_refill ? 1'h0 : _GEN_112; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  _GEN_121 = invalidate_refill ? 1'h0 : _GEN_113; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  _GEN_122 = invalidate_refill ? 1'h0 : _GEN_114; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  _GEN_123 = _T_9 ? _GEN_119 : sectored_entries_1_valid_0; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  _GEN_124 = _T_9 ? _GEN_120 : sectored_entries_1_valid_1; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  _GEN_125 = _T_9 ? _GEN_121 : sectored_entries_1_valid_2; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  _GEN_126 = _T_9 ? _GEN_122 : sectored_entries_1_valid_3; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  _T_11 = waddr == 3'h2; // @[TLB.scala 249:65]
  wire  _GEN_133 = _T_8 ? 1'h0 : sectored_entries_2_valid_0; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  _GEN_134 = _T_8 ? 1'h0 : sectored_entries_2_valid_1; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  _GEN_135 = _T_8 ? 1'h0 : sectored_entries_2_valid_2; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  _GEN_136 = _T_8 ? 1'h0 : sectored_entries_2_valid_3; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  _GEN_137 = (2'h0 == idx) | _GEN_133; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  _GEN_138 = (2'h1 == idx) | _GEN_134; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  _GEN_139 = (2'h2 == idx) | _GEN_135; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  _GEN_140 = (2'h3 == idx) | _GEN_136; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire [34:0] _GEN_141 = 2'h0 == idx ? _special_entry_data_0_T : sectored_entries_2_data_0; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] _GEN_142 = 2'h1 == idx ? _special_entry_data_0_T : sectored_entries_2_data_1; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] _GEN_143 = 2'h2 == idx ? _special_entry_data_0_T : sectored_entries_2_data_2; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] _GEN_144 = 2'h3 == idx ? _special_entry_data_0_T : sectored_entries_2_data_3; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire  _GEN_145 = invalidate_refill ? 1'h0 : _GEN_137; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  _GEN_146 = invalidate_refill ? 1'h0 : _GEN_138; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  _GEN_147 = invalidate_refill ? 1'h0 : _GEN_139; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  _GEN_148 = invalidate_refill ? 1'h0 : _GEN_140; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  _GEN_149 = _T_11 ? _GEN_145 : sectored_entries_2_valid_0; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  _GEN_150 = _T_11 ? _GEN_146 : sectored_entries_2_valid_1; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  _GEN_151 = _T_11 ? _GEN_147 : sectored_entries_2_valid_2; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  _GEN_152 = _T_11 ? _GEN_148 : sectored_entries_2_valid_3; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  _T_13 = waddr == 3'h3; // @[TLB.scala 249:65]
  wire  _GEN_159 = _T_8 ? 1'h0 : sectored_entries_3_valid_0; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  _GEN_160 = _T_8 ? 1'h0 : sectored_entries_3_valid_1; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  _GEN_161 = _T_8 ? 1'h0 : sectored_entries_3_valid_2; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  _GEN_162 = _T_8 ? 1'h0 : sectored_entries_3_valid_3; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  _GEN_163 = (2'h0 == idx) | _GEN_159; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  _GEN_164 = (2'h1 == idx) | _GEN_160; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  _GEN_165 = (2'h2 == idx) | _GEN_161; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  _GEN_166 = (2'h3 == idx) | _GEN_162; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire [34:0] _GEN_167 = 2'h0 == idx ? _special_entry_data_0_T : sectored_entries_3_data_0; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] _GEN_168 = 2'h1 == idx ? _special_entry_data_0_T : sectored_entries_3_data_1; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] _GEN_169 = 2'h2 == idx ? _special_entry_data_0_T : sectored_entries_3_data_2; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] _GEN_170 = 2'h3 == idx ? _special_entry_data_0_T : sectored_entries_3_data_3; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire  _GEN_171 = invalidate_refill ? 1'h0 : _GEN_163; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  _GEN_172 = invalidate_refill ? 1'h0 : _GEN_164; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  _GEN_173 = invalidate_refill ? 1'h0 : _GEN_165; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  _GEN_174 = invalidate_refill ? 1'h0 : _GEN_166; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  _GEN_175 = _T_13 ? _GEN_171 : sectored_entries_3_valid_0; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  _GEN_176 = _T_13 ? _GEN_172 : sectored_entries_3_valid_1; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  _GEN_177 = _T_13 ? _GEN_173 : sectored_entries_3_valid_2; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  _GEN_178 = _T_13 ? _GEN_174 : sectored_entries_3_valid_3; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  _T_15 = waddr == 3'h4; // @[TLB.scala 249:65]
  wire  _GEN_185 = _T_8 ? 1'h0 : sectored_entries_4_valid_0; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  _GEN_186 = _T_8 ? 1'h0 : sectored_entries_4_valid_1; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  _GEN_187 = _T_8 ? 1'h0 : sectored_entries_4_valid_2; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  _GEN_188 = _T_8 ? 1'h0 : sectored_entries_4_valid_3; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  _GEN_189 = (2'h0 == idx) | _GEN_185; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  _GEN_190 = (2'h1 == idx) | _GEN_186; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  _GEN_191 = (2'h2 == idx) | _GEN_187; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  _GEN_192 = (2'h3 == idx) | _GEN_188; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire [34:0] _GEN_193 = 2'h0 == idx ? _special_entry_data_0_T : sectored_entries_4_data_0; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] _GEN_194 = 2'h1 == idx ? _special_entry_data_0_T : sectored_entries_4_data_1; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] _GEN_195 = 2'h2 == idx ? _special_entry_data_0_T : sectored_entries_4_data_2; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] _GEN_196 = 2'h3 == idx ? _special_entry_data_0_T : sectored_entries_4_data_3; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire  _GEN_197 = invalidate_refill ? 1'h0 : _GEN_189; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  _GEN_198 = invalidate_refill ? 1'h0 : _GEN_190; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  _GEN_199 = invalidate_refill ? 1'h0 : _GEN_191; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  _GEN_200 = invalidate_refill ? 1'h0 : _GEN_192; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  _GEN_201 = _T_15 ? _GEN_197 : sectored_entries_4_valid_0; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  _GEN_202 = _T_15 ? _GEN_198 : sectored_entries_4_valid_1; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  _GEN_203 = _T_15 ? _GEN_199 : sectored_entries_4_valid_2; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  _GEN_204 = _T_15 ? _GEN_200 : sectored_entries_4_valid_3; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  _T_17 = waddr == 3'h5; // @[TLB.scala 249:65]
  wire  _GEN_211 = _T_8 ? 1'h0 : sectored_entries_5_valid_0; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  _GEN_212 = _T_8 ? 1'h0 : sectored_entries_5_valid_1; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  _GEN_213 = _T_8 ? 1'h0 : sectored_entries_5_valid_2; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  _GEN_214 = _T_8 ? 1'h0 : sectored_entries_5_valid_3; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  _GEN_215 = (2'h0 == idx) | _GEN_211; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  _GEN_216 = (2'h1 == idx) | _GEN_212; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  _GEN_217 = (2'h2 == idx) | _GEN_213; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  _GEN_218 = (2'h3 == idx) | _GEN_214; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire [34:0] _GEN_219 = 2'h0 == idx ? _special_entry_data_0_T : sectored_entries_5_data_0; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] _GEN_220 = 2'h1 == idx ? _special_entry_data_0_T : sectored_entries_5_data_1; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] _GEN_221 = 2'h2 == idx ? _special_entry_data_0_T : sectored_entries_5_data_2; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] _GEN_222 = 2'h3 == idx ? _special_entry_data_0_T : sectored_entries_5_data_3; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire  _GEN_223 = invalidate_refill ? 1'h0 : _GEN_215; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  _GEN_224 = invalidate_refill ? 1'h0 : _GEN_216; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  _GEN_225 = invalidate_refill ? 1'h0 : _GEN_217; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  _GEN_226 = invalidate_refill ? 1'h0 : _GEN_218; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  _GEN_227 = _T_17 ? _GEN_223 : sectored_entries_5_valid_0; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  _GEN_228 = _T_17 ? _GEN_224 : sectored_entries_5_valid_1; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  _GEN_229 = _T_17 ? _GEN_225 : sectored_entries_5_valid_2; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  _GEN_230 = _T_17 ? _GEN_226 : sectored_entries_5_valid_3; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  _T_19 = waddr == 3'h6; // @[TLB.scala 249:65]
  wire  _GEN_237 = _T_8 ? 1'h0 : sectored_entries_6_valid_0; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  _GEN_238 = _T_8 ? 1'h0 : sectored_entries_6_valid_1; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  _GEN_239 = _T_8 ? 1'h0 : sectored_entries_6_valid_2; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  _GEN_240 = _T_8 ? 1'h0 : sectored_entries_6_valid_3; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  _GEN_241 = (2'h0 == idx) | _GEN_237; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  _GEN_242 = (2'h1 == idx) | _GEN_238; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  _GEN_243 = (2'h2 == idx) | _GEN_239; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  _GEN_244 = (2'h3 == idx) | _GEN_240; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire [34:0] _GEN_245 = 2'h0 == idx ? _special_entry_data_0_T : sectored_entries_6_data_0; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] _GEN_246 = 2'h1 == idx ? _special_entry_data_0_T : sectored_entries_6_data_1; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] _GEN_247 = 2'h2 == idx ? _special_entry_data_0_T : sectored_entries_6_data_2; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] _GEN_248 = 2'h3 == idx ? _special_entry_data_0_T : sectored_entries_6_data_3; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire  _GEN_249 = invalidate_refill ? 1'h0 : _GEN_241; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  _GEN_250 = invalidate_refill ? 1'h0 : _GEN_242; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  _GEN_251 = invalidate_refill ? 1'h0 : _GEN_243; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  _GEN_252 = invalidate_refill ? 1'h0 : _GEN_244; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  _GEN_253 = _T_19 ? _GEN_249 : sectored_entries_6_valid_0; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  _GEN_254 = _T_19 ? _GEN_250 : sectored_entries_6_valid_1; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  _GEN_255 = _T_19 ? _GEN_251 : sectored_entries_6_valid_2; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  _GEN_256 = _T_19 ? _GEN_252 : sectored_entries_6_valid_3; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  _T_21 = waddr == 3'h7; // @[TLB.scala 249:65]
  wire  _GEN_263 = _T_8 ? 1'h0 : sectored_entries_7_valid_0; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  _GEN_264 = _T_8 ? 1'h0 : sectored_entries_7_valid_1; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  _GEN_265 = _T_8 ? 1'h0 : sectored_entries_7_valid_2; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  _GEN_266 = _T_8 ? 1'h0 : sectored_entries_7_valid_3; // @[TLB.scala 250:32 TLB.scala 126:38 TLB.scala 162:29]
  wire  _GEN_267 = (2'h0 == idx) | _GEN_263; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  _GEN_268 = (2'h1 == idx) | _GEN_264; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  _GEN_269 = (2'h2 == idx) | _GEN_265; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire  _GEN_270 = (2'h3 == idx) | _GEN_266; // @[TLB.scala 122:16 TLB.scala 122:16]
  wire [34:0] _GEN_271 = 2'h0 == idx ? _special_entry_data_0_T : sectored_entries_7_data_0; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] _GEN_272 = 2'h1 == idx ? _special_entry_data_0_T : sectored_entries_7_data_1; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] _GEN_273 = 2'h2 == idx ? _special_entry_data_0_T : sectored_entries_7_data_2; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire [34:0] _GEN_274 = 2'h3 == idx ? _special_entry_data_0_T : sectored_entries_7_data_3; // @[TLB.scala 123:15 TLB.scala 123:15 TLB.scala 162:29]
  wire  _GEN_275 = invalidate_refill ? 1'h0 : _GEN_267; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  _GEN_276 = invalidate_refill ? 1'h0 : _GEN_268; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  _GEN_277 = invalidate_refill ? 1'h0 : _GEN_269; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  _GEN_278 = invalidate_refill ? 1'h0 : _GEN_270; // @[TLB.scala 252:34 TLB.scala 126:38]
  wire  _GEN_279 = _T_21 ? _GEN_275 : sectored_entries_7_valid_0; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  _GEN_280 = _T_21 ? _GEN_276 : sectored_entries_7_valid_1; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  _GEN_281 = _T_21 ? _GEN_277 : sectored_entries_7_valid_2; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  _GEN_282 = _T_21 ? _GEN_278 : sectored_entries_7_valid_3; // @[TLB.scala 249:72 TLB.scala 162:29]
  wire  _GEN_291 = _T_2 ? _GEN_67 : superpage_entries_0_valid_0; // @[TLB.scala 242:54 TLB.scala 163:30]
  wire  _GEN_295 = _T_2 ? _GEN_71 : superpage_entries_1_valid_0; // @[TLB.scala 242:54 TLB.scala 163:30]
  wire  _GEN_299 = _T_2 ? _GEN_75 : superpage_entries_2_valid_0; // @[TLB.scala 242:54 TLB.scala 163:30]
  wire  _GEN_303 = _T_2 ? _GEN_79 : superpage_entries_3_valid_0; // @[TLB.scala 242:54 TLB.scala 163:30]
  wire  _GEN_305 = _T_2 ? sectored_entries_0_valid_0 : _GEN_97; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  _GEN_306 = _T_2 ? sectored_entries_0_valid_1 : _GEN_98; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  _GEN_307 = _T_2 ? sectored_entries_0_valid_2 : _GEN_99; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  _GEN_308 = _T_2 ? sectored_entries_0_valid_3 : _GEN_100; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  _GEN_315 = _T_2 ? sectored_entries_1_valid_0 : _GEN_123; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  _GEN_316 = _T_2 ? sectored_entries_1_valid_1 : _GEN_124; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  _GEN_317 = _T_2 ? sectored_entries_1_valid_2 : _GEN_125; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  _GEN_318 = _T_2 ? sectored_entries_1_valid_3 : _GEN_126; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  _GEN_325 = _T_2 ? sectored_entries_2_valid_0 : _GEN_149; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  _GEN_326 = _T_2 ? sectored_entries_2_valid_1 : _GEN_150; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  _GEN_327 = _T_2 ? sectored_entries_2_valid_2 : _GEN_151; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  _GEN_328 = _T_2 ? sectored_entries_2_valid_3 : _GEN_152; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  _GEN_335 = _T_2 ? sectored_entries_3_valid_0 : _GEN_175; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  _GEN_336 = _T_2 ? sectored_entries_3_valid_1 : _GEN_176; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  _GEN_337 = _T_2 ? sectored_entries_3_valid_2 : _GEN_177; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  _GEN_338 = _T_2 ? sectored_entries_3_valid_3 : _GEN_178; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  _GEN_345 = _T_2 ? sectored_entries_4_valid_0 : _GEN_201; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  _GEN_346 = _T_2 ? sectored_entries_4_valid_1 : _GEN_202; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  _GEN_347 = _T_2 ? sectored_entries_4_valid_2 : _GEN_203; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  _GEN_348 = _T_2 ? sectored_entries_4_valid_3 : _GEN_204; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  _GEN_355 = _T_2 ? sectored_entries_5_valid_0 : _GEN_227; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  _GEN_356 = _T_2 ? sectored_entries_5_valid_1 : _GEN_228; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  _GEN_357 = _T_2 ? sectored_entries_5_valid_2 : _GEN_229; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  _GEN_358 = _T_2 ? sectored_entries_5_valid_3 : _GEN_230; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  _GEN_365 = _T_2 ? sectored_entries_6_valid_0 : _GEN_253; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  _GEN_366 = _T_2 ? sectored_entries_6_valid_1 : _GEN_254; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  _GEN_367 = _T_2 ? sectored_entries_6_valid_2 : _GEN_255; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  _GEN_368 = _T_2 ? sectored_entries_6_valid_3 : _GEN_256; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  _GEN_375 = _T_2 ? sectored_entries_7_valid_0 : _GEN_279; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  _GEN_376 = _T_2 ? sectored_entries_7_valid_1 : _GEN_280; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  _GEN_377 = _T_2 ? sectored_entries_7_valid_2 : _GEN_281; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  _GEN_378 = _T_2 ? sectored_entries_7_valid_3 : _GEN_282; // @[TLB.scala 242:54 TLB.scala 162:29]
  wire  _GEN_387 = _T ? _GEN_64 : special_entry_valid_0; // @[TLB.scala 237:68 TLB.scala 164:56]
  wire  _GEN_391 = _T ? superpage_entries_0_valid_0 : _GEN_291; // @[TLB.scala 237:68 TLB.scala 163:30]
  wire  _GEN_395 = _T ? superpage_entries_1_valid_0 : _GEN_295; // @[TLB.scala 237:68 TLB.scala 163:30]
  wire  _GEN_399 = _T ? superpage_entries_2_valid_0 : _GEN_299; // @[TLB.scala 237:68 TLB.scala 163:30]
  wire  _GEN_403 = _T ? superpage_entries_3_valid_0 : _GEN_303; // @[TLB.scala 237:68 TLB.scala 163:30]
  wire  _GEN_405 = _T ? sectored_entries_0_valid_0 : _GEN_305; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  _GEN_406 = _T ? sectored_entries_0_valid_1 : _GEN_306; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  _GEN_407 = _T ? sectored_entries_0_valid_2 : _GEN_307; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  _GEN_408 = _T ? sectored_entries_0_valid_3 : _GEN_308; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  _GEN_415 = _T ? sectored_entries_1_valid_0 : _GEN_315; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  _GEN_416 = _T ? sectored_entries_1_valid_1 : _GEN_316; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  _GEN_417 = _T ? sectored_entries_1_valid_2 : _GEN_317; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  _GEN_418 = _T ? sectored_entries_1_valid_3 : _GEN_318; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  _GEN_425 = _T ? sectored_entries_2_valid_0 : _GEN_325; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  _GEN_426 = _T ? sectored_entries_2_valid_1 : _GEN_326; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  _GEN_427 = _T ? sectored_entries_2_valid_2 : _GEN_327; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  _GEN_428 = _T ? sectored_entries_2_valid_3 : _GEN_328; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  _GEN_435 = _T ? sectored_entries_3_valid_0 : _GEN_335; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  _GEN_436 = _T ? sectored_entries_3_valid_1 : _GEN_336; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  _GEN_437 = _T ? sectored_entries_3_valid_2 : _GEN_337; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  _GEN_438 = _T ? sectored_entries_3_valid_3 : _GEN_338; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  _GEN_445 = _T ? sectored_entries_4_valid_0 : _GEN_345; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  _GEN_446 = _T ? sectored_entries_4_valid_1 : _GEN_346; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  _GEN_447 = _T ? sectored_entries_4_valid_2 : _GEN_347; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  _GEN_448 = _T ? sectored_entries_4_valid_3 : _GEN_348; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  _GEN_455 = _T ? sectored_entries_5_valid_0 : _GEN_355; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  _GEN_456 = _T ? sectored_entries_5_valid_1 : _GEN_356; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  _GEN_457 = _T ? sectored_entries_5_valid_2 : _GEN_357; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  _GEN_458 = _T ? sectored_entries_5_valid_3 : _GEN_358; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  _GEN_465 = _T ? sectored_entries_6_valid_0 : _GEN_365; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  _GEN_466 = _T ? sectored_entries_6_valid_1 : _GEN_366; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  _GEN_467 = _T ? sectored_entries_6_valid_2 : _GEN_367; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  _GEN_468 = _T ? sectored_entries_6_valid_3 : _GEN_368; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  _GEN_475 = _T ? sectored_entries_7_valid_0 : _GEN_375; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  _GEN_476 = _T ? sectored_entries_7_valid_1 : _GEN_376; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  _GEN_477 = _T ? sectored_entries_7_valid_2 : _GEN_377; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  _GEN_478 = _T ? sectored_entries_7_valid_3 : _GEN_378; // @[TLB.scala 237:68 TLB.scala 162:29]
  wire  _GEN_487 = io_ptw_resp_valid ? _GEN_387 : special_entry_valid_0; // @[TLB.scala 217:20 TLB.scala 164:56]
  wire  _GEN_491 = io_ptw_resp_valid ? _GEN_391 : superpage_entries_0_valid_0; // @[TLB.scala 217:20 TLB.scala 163:30]
  wire  _GEN_495 = io_ptw_resp_valid ? _GEN_395 : superpage_entries_1_valid_0; // @[TLB.scala 217:20 TLB.scala 163:30]
  wire  _GEN_499 = io_ptw_resp_valid ? _GEN_399 : superpage_entries_2_valid_0; // @[TLB.scala 217:20 TLB.scala 163:30]
  wire  _GEN_503 = io_ptw_resp_valid ? _GEN_403 : superpage_entries_3_valid_0; // @[TLB.scala 217:20 TLB.scala 163:30]
  wire  _GEN_505 = io_ptw_resp_valid ? _GEN_405 : sectored_entries_0_valid_0; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  _GEN_506 = io_ptw_resp_valid ? _GEN_406 : sectored_entries_0_valid_1; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  _GEN_507 = io_ptw_resp_valid ? _GEN_407 : sectored_entries_0_valid_2; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  _GEN_508 = io_ptw_resp_valid ? _GEN_408 : sectored_entries_0_valid_3; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  _GEN_515 = io_ptw_resp_valid ? _GEN_415 : sectored_entries_1_valid_0; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  _GEN_516 = io_ptw_resp_valid ? _GEN_416 : sectored_entries_1_valid_1; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  _GEN_517 = io_ptw_resp_valid ? _GEN_417 : sectored_entries_1_valid_2; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  _GEN_518 = io_ptw_resp_valid ? _GEN_418 : sectored_entries_1_valid_3; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  _GEN_525 = io_ptw_resp_valid ? _GEN_425 : sectored_entries_2_valid_0; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  _GEN_526 = io_ptw_resp_valid ? _GEN_426 : sectored_entries_2_valid_1; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  _GEN_527 = io_ptw_resp_valid ? _GEN_427 : sectored_entries_2_valid_2; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  _GEN_528 = io_ptw_resp_valid ? _GEN_428 : sectored_entries_2_valid_3; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  _GEN_535 = io_ptw_resp_valid ? _GEN_435 : sectored_entries_3_valid_0; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  _GEN_536 = io_ptw_resp_valid ? _GEN_436 : sectored_entries_3_valid_1; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  _GEN_537 = io_ptw_resp_valid ? _GEN_437 : sectored_entries_3_valid_2; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  _GEN_538 = io_ptw_resp_valid ? _GEN_438 : sectored_entries_3_valid_3; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  _GEN_545 = io_ptw_resp_valid ? _GEN_445 : sectored_entries_4_valid_0; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  _GEN_546 = io_ptw_resp_valid ? _GEN_446 : sectored_entries_4_valid_1; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  _GEN_547 = io_ptw_resp_valid ? _GEN_447 : sectored_entries_4_valid_2; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  _GEN_548 = io_ptw_resp_valid ? _GEN_448 : sectored_entries_4_valid_3; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  _GEN_555 = io_ptw_resp_valid ? _GEN_455 : sectored_entries_5_valid_0; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  _GEN_556 = io_ptw_resp_valid ? _GEN_456 : sectored_entries_5_valid_1; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  _GEN_557 = io_ptw_resp_valid ? _GEN_457 : sectored_entries_5_valid_2; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  _GEN_558 = io_ptw_resp_valid ? _GEN_458 : sectored_entries_5_valid_3; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  _GEN_565 = io_ptw_resp_valid ? _GEN_465 : sectored_entries_6_valid_0; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  _GEN_566 = io_ptw_resp_valid ? _GEN_466 : sectored_entries_6_valid_1; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  _GEN_567 = io_ptw_resp_valid ? _GEN_467 : sectored_entries_6_valid_2; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  _GEN_568 = io_ptw_resp_valid ? _GEN_468 : sectored_entries_6_valid_3; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  _GEN_575 = io_ptw_resp_valid ? _GEN_475 : sectored_entries_7_valid_0; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  _GEN_576 = io_ptw_resp_valid ? _GEN_476 : sectored_entries_7_valid_1; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  _GEN_577 = io_ptw_resp_valid ? _GEN_477 : sectored_entries_7_valid_2; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire  _GEN_578 = io_ptw_resp_valid ? _GEN_478 : sectored_entries_7_valid_3; // @[TLB.scala 217:20 TLB.scala 162:29]
  wire [5:0] ptw_ae_array_left = {entries_barrier_5_io_y_ae,entries_barrier_4_io_y_ae,entries_barrier_3_io_y_ae,
    entries_barrier_2_io_y_ae,entries_barrier_1_io_y_ae,entries_barrier_io_y_ae}; // @[Cat.scala 29:58]
  wire [13:0] ptw_ae_array = {1'h0,entries_barrier_12_io_y_ae,entries_barrier_11_io_y_ae,entries_barrier_10_io_y_ae,
    entries_barrier_9_io_y_ae,entries_barrier_8_io_y_ae,entries_barrier_7_io_y_ae,entries_barrier_6_io_y_ae,
    ptw_ae_array_left}; // @[Cat.scala 29:58]
  wire [5:0] priv_rw_ok_left = {entries_barrier_5_io_y_u,entries_barrier_4_io_y_u,entries_barrier_3_io_y_u,
    entries_barrier_2_io_y_u,entries_barrier_1_io_y_u,entries_barrier_io_y_u}; // @[Cat.scala 29:58]
  wire [12:0] _priv_rw_ok_T_2 = {entries_barrier_12_io_y_u,entries_barrier_11_io_y_u,entries_barrier_10_io_y_u,
    entries_barrier_9_io_y_u,entries_barrier_8_io_y_u,entries_barrier_7_io_y_u,entries_barrier_6_io_y_u,priv_rw_ok_left}
    ; // @[Cat.scala 29:58]
  wire [12:0] _priv_rw_ok_T_5 = ~_priv_rw_ok_T_2; // @[TLB.scala 261:98]
  wire [12:0] priv_x_ok = priv_s ? _priv_rw_ok_T_5 : _priv_rw_ok_T_2; // @[TLB.scala 262:22]
  wire [5:0] r_array_left_1 = {entries_barrier_5_io_y_sx,entries_barrier_4_io_y_sx,entries_barrier_3_io_y_sx,
    entries_barrier_2_io_y_sx,entries_barrier_1_io_y_sx,entries_barrier_io_y_sx}; // @[Cat.scala 29:58]
  wire [12:0] _r_array_T_1 = {entries_barrier_12_io_y_sx,entries_barrier_11_io_y_sx,entries_barrier_10_io_y_sx,
    entries_barrier_9_io_y_sx,entries_barrier_8_io_y_sx,entries_barrier_7_io_y_sx,entries_barrier_6_io_y_sx,
    r_array_left_1}; // @[Cat.scala 29:58]
  wire [12:0] x_array_left_1 = priv_x_ok & _r_array_T_1; // @[TLB.scala 265:39]
  wire [13:0] x_array = {1'h1,x_array_left_1}; // @[Cat.scala 29:58]
  wire [13:0] _pr_array_T_2 = ~ptw_ae_array; // @[TLB.scala 266:89]
  wire [1:0] px_array_right = prot_x ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [5:0] px_array_left = {normal_entries_barrier_5_io_y_px,normal_entries_barrier_4_io_y_px,
    normal_entries_barrier_3_io_y_px,normal_entries_barrier_2_io_y_px,normal_entries_barrier_1_io_y_px,
    normal_entries_barrier_io_y_px}; // @[Cat.scala 29:58]
  wire [13:0] _px_array_T_1 = {px_array_right,normal_entries_barrier_11_io_y_px,normal_entries_barrier_10_io_y_px,
    normal_entries_barrier_9_io_y_px,normal_entries_barrier_8_io_y_px,normal_entries_barrier_7_io_y_px,
    normal_entries_barrier_6_io_y_px,px_array_left}; // @[Cat.scala 29:58]
  wire [13:0] px_array = _px_array_T_1 & _pr_array_T_2; // @[TLB.scala 268:87]
  wire [1:0] c_array_right = cacheable ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [5:0] c_array_left = {normal_entries_barrier_5_io_y_c,normal_entries_barrier_4_io_y_c,
    normal_entries_barrier_3_io_y_c,normal_entries_barrier_2_io_y_c,normal_entries_barrier_1_io_y_c,
    normal_entries_barrier_io_y_c}; // @[Cat.scala 29:58]
  wire [13:0] c_array = {c_array_right,normal_entries_barrier_11_io_y_c,normal_entries_barrier_10_io_y_c,
    normal_entries_barrier_9_io_y_c,normal_entries_barrier_8_io_y_c,normal_entries_barrier_7_io_y_c,
    normal_entries_barrier_6_io_y_c,c_array_left}; // @[Cat.scala 29:58]
  wire [39:0] bad_va_maskedVAddr = io_req_bits_vaddr & 40'hc000000000; // @[TLB.scala 285:43]
  wire  _bad_va_T_4 = ~((bad_va_maskedVAddr == 40'h0) | (bad_va_maskedVAddr == 40'hc000000000)); // @[TLB.scala 286:47]
  wire  bad_va = vm_enabled & _bad_va_T_4; // @[TLB.scala 280:117]
  wire [13:0] _pf_inst_array_T = x_array | ptw_ae_array; // @[TLB.scala 318:33]
  wire [13:0] pf_inst_array = ~_pf_inst_array_T; // @[TLB.scala 318:23]
  wire  tlb_hit = |real_hits; // @[TLB.scala 320:27]
  wire  tlb_miss = (vm_enabled & (~bad_va)) & (~tlb_hit); // @[TLB.scala 321:40]
  reg [6:0] state_reg; // @[Replacement.scala 158:30]
  reg [2:0] state_reg_1; // @[Replacement.scala 158:30]
  wire  _T_23 = io_req_valid & vm_enabled; // @[TLB.scala 325:22]
  wire  _T_30 = ((((((sector_hits_0 | sector_hits_1) | sector_hits_2) | sector_hits_3) | sector_hits_4) | sector_hits_5)
     | sector_hits_6) | sector_hits_7; // @[package.scala 64:59]
  wire [7:0] _T_31 = {sector_hits_7,sector_hits_6,sector_hits_5,sector_hits_4,sector_hits_3,sector_hits_2,sector_hits_1,
    sector_hits_0}; // @[Cat.scala 29:58]
  wire [3:0] hi = _T_31[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] lo = _T_31[3:0]; // @[OneHot.scala 31:18]
  wire  right_1 = |hi; // @[OneHot.scala 32:14]
  wire [3:0] _T_32 = hi | lo; // @[OneHot.scala 32:28]
  wire [1:0] hi_1 = _T_32[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] lo_1 = _T_32[1:0]; // @[OneHot.scala 31:18]
  wire  right_2 = |hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _T_33 = hi_1 | lo_1; // @[OneHot.scala 32:28]
  wire  left_1 = _T_33[1]; // @[CircuitMath.scala 30:8]
  wire [2:0] state_reg_touch_way_sized = {right_1,right_2,left_1}; // @[Cat.scala 29:58]
  wire  state_reg_right_right = ~(state_reg_touch_way_sized[2]); // @[Replacement.scala 186:33]
  wire [2:0] state_reg_left_subtree_state = state_reg[5:3]; // @[package.scala 143:13]
  wire [2:0] state_reg_right_subtree_state = state_reg[2:0]; // @[Replacement.scala 188:38]
  wire  state_reg_right_right_1 = ~(state_reg_touch_way_sized[1]); // @[Replacement.scala 186:33]
  wire  state_reg_left_subtree_state_1 = state_reg_left_subtree_state[1]; // @[package.scala 143:13]
  wire  state_reg_right_subtree_state_1 = state_reg_left_subtree_state[0]; // @[Replacement.scala 188:38]
  wire  _state_reg_T_3 = ~(state_reg_touch_way_sized[0]); // @[Replacement.scala 208:7]
  wire  state_reg_right_left = state_reg_right_right_1 ? state_reg_left_subtree_state_1 : _state_reg_T_3; // @[Replacement.scala 193:16]
  wire  state_reg_left = state_reg_right_right_1 ? _state_reg_T_3 : state_reg_right_subtree_state_1; // @[Replacement.scala 196:16]
  wire [2:0] _state_reg_T_7 = {state_reg_right_right_1,state_reg_right_left,state_reg_left}; // @[Cat.scala 29:58]
  wire [2:0] state_reg_right_left_1 = state_reg_right_right ? state_reg_left_subtree_state : _state_reg_T_7; // @[Replacement.scala 193:16]
  wire  state_reg_left_subtree_state_2 = state_reg_right_subtree_state[1]; // @[package.scala 143:13]
  wire  state_reg_right_subtree_state_2 = state_reg_right_subtree_state[0]; // @[Replacement.scala 188:38]
  wire  state_reg_right_left_2 = state_reg_right_right_1 ? state_reg_left_subtree_state_2 : _state_reg_T_3; // @[Replacement.scala 193:16]
  wire  state_reg_left_1 = state_reg_right_right_1 ? _state_reg_T_3 : state_reg_right_subtree_state_2; // @[Replacement.scala 196:16]
  wire [2:0] _state_reg_T_15 = {state_reg_right_right_1,state_reg_right_left_2,state_reg_left_1}; // @[Cat.scala 29:58]
  wire [2:0] state_reg_left_2 = state_reg_right_right ? _state_reg_T_15 : state_reg_right_subtree_state; // @[Replacement.scala 196:16]
  wire [6:0] _state_reg_T_16 = {state_reg_right_right,state_reg_right_left_1,state_reg_left_2}; // @[Cat.scala 29:58]
  wire  _T_37 = ((superpage_hits_0 | superpage_hits_1) | superpage_hits_2) | superpage_hits_3; // @[package.scala 64:59]
  wire [3:0] _T_38 = {superpage_hits_3,superpage_hits_2,superpage_hits_1,superpage_hits_0}; // @[Cat.scala 29:58]
  wire [1:0] hi_2 = _T_38[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] lo_2 = _T_38[1:0]; // @[OneHot.scala 31:18]
  wire  right_4 = |hi_2; // @[OneHot.scala 32:14]
  wire [1:0] _T_39 = hi_2 | lo_2; // @[OneHot.scala 32:28]
  wire  left_4 = _T_39[1]; // @[CircuitMath.scala 30:8]
  wire [1:0] state_reg_1_touch_way_sized = {right_4,left_4}; // @[Cat.scala 29:58]
  wire  state_reg_1_right_right = ~(state_reg_1_touch_way_sized[1]); // @[Replacement.scala 186:33]
  wire  state_reg_1_left_subtree_state = state_reg_1[1]; // @[package.scala 143:13]
  wire  state_reg_1_right_subtree_state = state_reg_1[0]; // @[Replacement.scala 188:38]
  wire  _state_reg_1_T_2 = ~(state_reg_1_touch_way_sized[0]); // @[Replacement.scala 208:7]
  wire  state_reg_1_right_left = state_reg_1_right_right ? state_reg_1_left_subtree_state : _state_reg_1_T_2; // @[Replacement.scala 193:16]
  wire  state_reg_1_left = state_reg_1_right_right ? _state_reg_1_T_2 : state_reg_1_right_subtree_state; // @[Replacement.scala 196:16]
  wire [2:0] _state_reg_1_T_6 = {state_reg_1_right_right,state_reg_1_right_left,state_reg_1_left}; // @[Cat.scala 29:58]
  wire  multipleHits_leftOne = real_hits[0]; // @[Misc.scala 180:37]
  wire  multipleHits_leftOne_1 = real_hits[1]; // @[Misc.scala 180:37]
  wire  multipleHits_rightOne = real_hits[2]; // @[Misc.scala 181:39]
  wire  multipleHits_rightOne_1 = multipleHits_leftOne_1 | multipleHits_rightOne; // @[Misc.scala 182:16]
  wire  multipleHits_rightTwo = multipleHits_leftOne_1 & multipleHits_rightOne; // @[Misc.scala 182:61]
  wire  multipleHits_leftOne_2 = multipleHits_leftOne | multipleHits_rightOne_1; // @[Misc.scala 182:16]
  wire  multipleHits_leftTwo = multipleHits_rightTwo | (multipleHits_leftOne & multipleHits_rightOne_1); // @[Misc.scala 182:49]
  wire  multipleHits_leftOne_3 = real_hits[3]; // @[Misc.scala 180:37]
  wire  multipleHits_leftOne_4 = real_hits[4]; // @[Misc.scala 180:37]
  wire  multipleHits_rightOne_2 = real_hits[5]; // @[Misc.scala 181:39]
  wire  multipleHits_rightOne_3 = multipleHits_leftOne_4 | multipleHits_rightOne_2; // @[Misc.scala 182:16]
  wire  multipleHits_rightTwo_1 = multipleHits_leftOne_4 & multipleHits_rightOne_2; // @[Misc.scala 182:61]
  wire  multipleHits_rightOne_4 = multipleHits_leftOne_3 | multipleHits_rightOne_3; // @[Misc.scala 182:16]
  wire  multipleHits_rightTwo_2 = multipleHits_rightTwo_1 | (multipleHits_leftOne_3 & multipleHits_rightOne_3); // @[Misc.scala 182:49]
  wire  multipleHits_leftOne_5 = multipleHits_leftOne_2 | multipleHits_rightOne_4; // @[Misc.scala 182:16]
  wire  multipleHits_leftTwo_1 = (multipleHits_leftTwo | multipleHits_rightTwo_2) | (multipleHits_leftOne_2 &
    multipleHits_rightOne_4); // @[Misc.scala 182:49]
  wire  multipleHits_leftOne_6 = real_hits[6]; // @[Misc.scala 180:37]
  wire  multipleHits_leftOne_7 = real_hits[7]; // @[Misc.scala 180:37]
  wire  multipleHits_rightOne_5 = real_hits[8]; // @[Misc.scala 181:39]
  wire  multipleHits_rightOne_6 = multipleHits_leftOne_7 | multipleHits_rightOne_5; // @[Misc.scala 182:16]
  wire  multipleHits_rightTwo_3 = multipleHits_leftOne_7 & multipleHits_rightOne_5; // @[Misc.scala 182:61]
  wire  multipleHits_leftOne_8 = multipleHits_leftOne_6 | multipleHits_rightOne_6; // @[Misc.scala 182:16]
  wire  multipleHits_leftTwo_2 = multipleHits_rightTwo_3 | (multipleHits_leftOne_6 & multipleHits_rightOne_6); // @[Misc.scala 182:49]
  wire  multipleHits_leftOne_9 = real_hits[9]; // @[Misc.scala 180:37]
  wire  multipleHits_rightOne_7 = real_hits[10]; // @[Misc.scala 181:39]
  wire  multipleHits_leftOne_10 = multipleHits_leftOne_9 | multipleHits_rightOne_7; // @[Misc.scala 182:16]
  wire  multipleHits_leftTwo_3 = multipleHits_leftOne_9 & multipleHits_rightOne_7; // @[Misc.scala 182:61]
  wire  multipleHits_leftOne_11 = real_hits[11]; // @[Misc.scala 180:37]
  wire  multipleHits_rightOne_8 = real_hits[12]; // @[Misc.scala 181:39]
  wire  multipleHits_rightOne_9 = multipleHits_leftOne_11 | multipleHits_rightOne_8; // @[Misc.scala 182:16]
  wire  multipleHits_rightTwo_4 = multipleHits_leftOne_11 & multipleHits_rightOne_8; // @[Misc.scala 182:61]
  wire  multipleHits_rightOne_10 = multipleHits_leftOne_10 | multipleHits_rightOne_9; // @[Misc.scala 182:16]
  wire  multipleHits_rightTwo_5 = (multipleHits_leftTwo_3 | multipleHits_rightTwo_4) | (multipleHits_leftOne_10 &
    multipleHits_rightOne_9); // @[Misc.scala 182:49]
  wire  multipleHits_rightOne_11 = multipleHits_leftOne_8 | multipleHits_rightOne_10; // @[Misc.scala 182:16]
  wire  multipleHits_rightTwo_6 = (multipleHits_leftTwo_2 | multipleHits_rightTwo_5) | (multipleHits_leftOne_8 &
    multipleHits_rightOne_10); // @[Misc.scala 182:49]
  wire  multipleHits = (multipleHits_leftTwo_1 | multipleHits_rightTwo_6) | (multipleHits_leftOne_5 &
    multipleHits_rightOne_11); // @[Misc.scala 182:49]
  wire [13:0] _io_resp_pf_inst_T = pf_inst_array & hits; // @[TLB.scala 340:47]
  wire [13:0] _io_resp_ae_inst_T = ~px_array; // @[TLB.scala 343:23]
  wire [13:0] _io_resp_ae_inst_T_1 = _io_resp_ae_inst_T & hits; // @[TLB.scala 343:33]
  wire [13:0] _io_resp_cacheable_T = c_array & hits; // @[TLB.scala 347:33]
  wire  _T_41 = io_req_ready & io_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_42 = _T_41 & tlb_miss; // @[TLB.scala 359:25]
  wire  r_superpage_repl_addr_right = state_reg_1[2]; // @[Replacement.scala 233:38]
  wire  r_superpage_repl_addr_left = r_superpage_repl_addr_right ? state_reg_1_left_subtree_state :
    state_reg_1_right_subtree_state; // @[Replacement.scala 240:16]
  wire [1:0] _r_superpage_repl_addr_T_2 = {r_superpage_repl_addr_right,r_superpage_repl_addr_left}; // @[Cat.scala 29:58]
  wire [3:0] r_superpage_repl_addr_valids = {superpage_entries_3_valid_0,superpage_entries_2_valid_0,
    superpage_entries_1_valid_0,superpage_entries_0_valid_0}; // @[Cat.scala 29:58]
  wire [3:0] _r_superpage_repl_addr_T_4 = ~r_superpage_repl_addr_valids; // @[TLB.scala 407:43]
  wire [1:0] _r_superpage_repl_addr_T_9 = _r_superpage_repl_addr_T_4[2] ? 2'h2 : 2'h3; // @[Mux.scala 47:69]
  wire  r_sectored_repl_addr_right = state_reg[6]; // @[Replacement.scala 233:38]
  wire  r_sectored_repl_addr_right_1 = state_reg_left_subtree_state[2]; // @[Replacement.scala 233:38]
  wire  r_sectored_repl_addr_left = r_sectored_repl_addr_right_1 ? state_reg_left_subtree_state_1 :
    state_reg_right_subtree_state_1; // @[Replacement.scala 240:16]
  wire [1:0] _r_sectored_repl_addr_T_2 = {r_sectored_repl_addr_right_1,r_sectored_repl_addr_left}; // @[Cat.scala 29:58]
  wire  r_sectored_repl_addr_right_2 = state_reg_right_subtree_state[2]; // @[Replacement.scala 233:38]
  wire  r_sectored_repl_addr_left_1 = r_sectored_repl_addr_right_2 ? state_reg_left_subtree_state_2 :
    state_reg_right_subtree_state_2; // @[Replacement.scala 240:16]
  wire [1:0] _r_sectored_repl_addr_T_5 = {r_sectored_repl_addr_right_2,r_sectored_repl_addr_left_1}; // @[Cat.scala 29:58]
  wire [1:0] r_sectored_repl_addr_left_2 = r_sectored_repl_addr_right ? _r_sectored_repl_addr_T_2 :
    _r_sectored_repl_addr_T_5; // @[Replacement.scala 240:16]
  wire [2:0] _r_sectored_repl_addr_T_6 = {r_sectored_repl_addr_right,r_sectored_repl_addr_left_2}; // @[Cat.scala 29:58]
  wire [7:0] r_sectored_repl_addr_valids = {_sector_hits_T_44,_sector_hits_T_38,_sector_hits_T_32,_sector_hits_T_26,
    _sector_hits_T_20,_sector_hits_T_14,_sector_hits_T_8,_sector_hits_T_2}; // @[Cat.scala 29:58]
  wire [7:0] _r_sectored_repl_addr_T_8 = ~r_sectored_repl_addr_valids; // @[TLB.scala 407:43]
  wire [2:0] _r_sectored_repl_addr_T_17 = _r_sectored_repl_addr_T_8[6] ? 3'h6 : 3'h7; // @[Mux.scala 47:69]
  wire [2:0] _r_sectored_repl_addr_T_18 = _r_sectored_repl_addr_T_8[5] ? 3'h5 : _r_sectored_repl_addr_T_17; // @[Mux.scala 47:69]
  wire [2:0] _r_sectored_repl_addr_T_19 = _r_sectored_repl_addr_T_8[4] ? 3'h4 : _r_sectored_repl_addr_T_18; // @[Mux.scala 47:69]
  wire [2:0] _r_sectored_repl_addr_T_20 = _r_sectored_repl_addr_T_8[3] ? 3'h3 : _r_sectored_repl_addr_T_19; // @[Mux.scala 47:69]
  wire [2:0] _r_sectored_repl_addr_T_21 = _r_sectored_repl_addr_T_8[2] ? 3'h2 : _r_sectored_repl_addr_T_20; // @[Mux.scala 47:69]
  wire [1:0] _GEN_653 = _T_42 ? 2'h1 : state; // @[TLB.scala 359:38 TLB.scala 360:13 TLB.scala 169:18]
  wire [1:0] _GEN_659 = io_sfence_valid ? 2'h0 : _GEN_653; // @[TLB.scala 369:21 TLB.scala 369:29]
  wire [1:0] _state_T = io_sfence_valid ? 2'h3 : 2'h2; // @[TLB.scala 370:45]
  wire [1:0] _GEN_660 = io_ptw_req_ready ? _state_T : _GEN_659; // @[TLB.scala 370:31 TLB.scala 370:39]
  wire [1:0] _GEN_661 = io_kill ? 2'h0 : _GEN_660; // @[TLB.scala 371:22 TLB.scala 371:30]
  wire  _T_45 = (state == 2'h2) & io_sfence_valid; // @[TLB.scala 373:28]
  wire  _GEN_665 = 2'h0 == hitsVec_idx ? 1'h0 : _GEN_505; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  _GEN_666 = 2'h1 == hitsVec_idx ? 1'h0 : _GEN_506; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  _GEN_667 = 2'h2 == hitsVec_idx ? 1'h0 : _GEN_507; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  _GEN_668 = 2'h3 == hitsVec_idx ? 1'h0 : _GEN_508; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  _GEN_669 = _sector_hits_T_5 ? _GEN_665 : _GEN_505; // @[TLB.scala 131:34]
  wire  _GEN_670 = _sector_hits_T_5 ? _GEN_666 : _GEN_506; // @[TLB.scala 131:34]
  wire  _GEN_671 = _sector_hits_T_5 ? _GEN_667 : _GEN_507; // @[TLB.scala 131:34]
  wire  _GEN_672 = _sector_hits_T_5 ? _GEN_668 : _GEN_508; // @[TLB.scala 131:34]
  wire  _T_59 = (_sector_hits_T_3[26:18]) == 9'h0; // @[TLB.scala 135:61]
  wire  _GEN_673 = sectored_entries_0_data_0[0] ? 1'h0 : _GEN_669; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  _GEN_674 = sectored_entries_0_data_1[0] ? 1'h0 : _GEN_670; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  _GEN_675 = sectored_entries_0_data_2[0] ? 1'h0 : _GEN_671; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  _GEN_676 = sectored_entries_0_data_3[0] ? 1'h0 : _GEN_672; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  _T_188 = ~(sectored_entries_0_data_0[13]); // @[TLB.scala 143:13]
  wire  _GEN_681 = _T_188 ? 1'h0 : _GEN_505; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _T_189 = ~(sectored_entries_0_data_1[13]); // @[TLB.scala 143:13]
  wire  _GEN_682 = _T_189 ? 1'h0 : _GEN_506; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _T_190 = ~(sectored_entries_0_data_2[13]); // @[TLB.scala 143:13]
  wire  _GEN_683 = _T_190 ? 1'h0 : _GEN_507; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _T_191 = ~(sectored_entries_0_data_3[13]); // @[TLB.scala 143:13]
  wire  _GEN_684 = _T_191 ? 1'h0 : _GEN_508; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _GEN_685 = io_sfence_bits_rs2 & _GEN_681; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _GEN_686 = io_sfence_bits_rs2 & _GEN_682; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _GEN_687 = io_sfence_bits_rs2 & _GEN_683; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _GEN_688 = io_sfence_bits_rs2 & _GEN_684; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _GEN_693 = 2'h0 == hitsVec_idx ? 1'h0 : _GEN_515; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  _GEN_694 = 2'h1 == hitsVec_idx ? 1'h0 : _GEN_516; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  _GEN_695 = 2'h2 == hitsVec_idx ? 1'h0 : _GEN_517; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  _GEN_696 = 2'h3 == hitsVec_idx ? 1'h0 : _GEN_518; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  _GEN_697 = _sector_hits_T_11 ? _GEN_693 : _GEN_515; // @[TLB.scala 131:34]
  wire  _GEN_698 = _sector_hits_T_11 ? _GEN_694 : _GEN_516; // @[TLB.scala 131:34]
  wire  _GEN_699 = _sector_hits_T_11 ? _GEN_695 : _GEN_517; // @[TLB.scala 131:34]
  wire  _GEN_700 = _sector_hits_T_11 ? _GEN_696 : _GEN_518; // @[TLB.scala 131:34]
  wire  _T_198 = (_sector_hits_T_9[26:18]) == 9'h0; // @[TLB.scala 135:61]
  wire  _GEN_701 = sectored_entries_1_data_0[0] ? 1'h0 : _GEN_697; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  _GEN_702 = sectored_entries_1_data_1[0] ? 1'h0 : _GEN_698; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  _GEN_703 = sectored_entries_1_data_2[0] ? 1'h0 : _GEN_699; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  _GEN_704 = sectored_entries_1_data_3[0] ? 1'h0 : _GEN_700; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  _T_327 = ~(sectored_entries_1_data_0[13]); // @[TLB.scala 143:13]
  wire  _GEN_709 = _T_327 ? 1'h0 : _GEN_515; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _T_328 = ~(sectored_entries_1_data_1[13]); // @[TLB.scala 143:13]
  wire  _GEN_710 = _T_328 ? 1'h0 : _GEN_516; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _T_329 = ~(sectored_entries_1_data_2[13]); // @[TLB.scala 143:13]
  wire  _GEN_711 = _T_329 ? 1'h0 : _GEN_517; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _T_330 = ~(sectored_entries_1_data_3[13]); // @[TLB.scala 143:13]
  wire  _GEN_712 = _T_330 ? 1'h0 : _GEN_518; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _GEN_713 = io_sfence_bits_rs2 & _GEN_709; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _GEN_714 = io_sfence_bits_rs2 & _GEN_710; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _GEN_715 = io_sfence_bits_rs2 & _GEN_711; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _GEN_716 = io_sfence_bits_rs2 & _GEN_712; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _GEN_721 = 2'h0 == hitsVec_idx ? 1'h0 : _GEN_525; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  _GEN_722 = 2'h1 == hitsVec_idx ? 1'h0 : _GEN_526; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  _GEN_723 = 2'h2 == hitsVec_idx ? 1'h0 : _GEN_527; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  _GEN_724 = 2'h3 == hitsVec_idx ? 1'h0 : _GEN_528; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  _GEN_725 = _sector_hits_T_17 ? _GEN_721 : _GEN_525; // @[TLB.scala 131:34]
  wire  _GEN_726 = _sector_hits_T_17 ? _GEN_722 : _GEN_526; // @[TLB.scala 131:34]
  wire  _GEN_727 = _sector_hits_T_17 ? _GEN_723 : _GEN_527; // @[TLB.scala 131:34]
  wire  _GEN_728 = _sector_hits_T_17 ? _GEN_724 : _GEN_528; // @[TLB.scala 131:34]
  wire  _T_337 = (_sector_hits_T_15[26:18]) == 9'h0; // @[TLB.scala 135:61]
  wire  _GEN_729 = sectored_entries_2_data_0[0] ? 1'h0 : _GEN_725; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  _GEN_730 = sectored_entries_2_data_1[0] ? 1'h0 : _GEN_726; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  _GEN_731 = sectored_entries_2_data_2[0] ? 1'h0 : _GEN_727; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  _GEN_732 = sectored_entries_2_data_3[0] ? 1'h0 : _GEN_728; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  _T_466 = ~(sectored_entries_2_data_0[13]); // @[TLB.scala 143:13]
  wire  _GEN_737 = _T_466 ? 1'h0 : _GEN_525; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _T_467 = ~(sectored_entries_2_data_1[13]); // @[TLB.scala 143:13]
  wire  _GEN_738 = _T_467 ? 1'h0 : _GEN_526; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _T_468 = ~(sectored_entries_2_data_2[13]); // @[TLB.scala 143:13]
  wire  _GEN_739 = _T_468 ? 1'h0 : _GEN_527; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _T_469 = ~(sectored_entries_2_data_3[13]); // @[TLB.scala 143:13]
  wire  _GEN_740 = _T_469 ? 1'h0 : _GEN_528; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _GEN_741 = io_sfence_bits_rs2 & _GEN_737; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _GEN_742 = io_sfence_bits_rs2 & _GEN_738; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _GEN_743 = io_sfence_bits_rs2 & _GEN_739; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _GEN_744 = io_sfence_bits_rs2 & _GEN_740; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _GEN_749 = 2'h0 == hitsVec_idx ? 1'h0 : _GEN_535; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  _GEN_750 = 2'h1 == hitsVec_idx ? 1'h0 : _GEN_536; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  _GEN_751 = 2'h2 == hitsVec_idx ? 1'h0 : _GEN_537; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  _GEN_752 = 2'h3 == hitsVec_idx ? 1'h0 : _GEN_538; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  _GEN_753 = _sector_hits_T_23 ? _GEN_749 : _GEN_535; // @[TLB.scala 131:34]
  wire  _GEN_754 = _sector_hits_T_23 ? _GEN_750 : _GEN_536; // @[TLB.scala 131:34]
  wire  _GEN_755 = _sector_hits_T_23 ? _GEN_751 : _GEN_537; // @[TLB.scala 131:34]
  wire  _GEN_756 = _sector_hits_T_23 ? _GEN_752 : _GEN_538; // @[TLB.scala 131:34]
  wire  _T_476 = (_sector_hits_T_21[26:18]) == 9'h0; // @[TLB.scala 135:61]
  wire  _GEN_757 = sectored_entries_3_data_0[0] ? 1'h0 : _GEN_753; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  _GEN_758 = sectored_entries_3_data_1[0] ? 1'h0 : _GEN_754; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  _GEN_759 = sectored_entries_3_data_2[0] ? 1'h0 : _GEN_755; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  _GEN_760 = sectored_entries_3_data_3[0] ? 1'h0 : _GEN_756; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  _T_605 = ~(sectored_entries_3_data_0[13]); // @[TLB.scala 143:13]
  wire  _GEN_765 = _T_605 ? 1'h0 : _GEN_535; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _T_606 = ~(sectored_entries_3_data_1[13]); // @[TLB.scala 143:13]
  wire  _GEN_766 = _T_606 ? 1'h0 : _GEN_536; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _T_607 = ~(sectored_entries_3_data_2[13]); // @[TLB.scala 143:13]
  wire  _GEN_767 = _T_607 ? 1'h0 : _GEN_537; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _T_608 = ~(sectored_entries_3_data_3[13]); // @[TLB.scala 143:13]
  wire  _GEN_768 = _T_608 ? 1'h0 : _GEN_538; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _GEN_769 = io_sfence_bits_rs2 & _GEN_765; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _GEN_770 = io_sfence_bits_rs2 & _GEN_766; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _GEN_771 = io_sfence_bits_rs2 & _GEN_767; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _GEN_772 = io_sfence_bits_rs2 & _GEN_768; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _GEN_777 = 2'h0 == hitsVec_idx ? 1'h0 : _GEN_545; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  _GEN_778 = 2'h1 == hitsVec_idx ? 1'h0 : _GEN_546; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  _GEN_779 = 2'h2 == hitsVec_idx ? 1'h0 : _GEN_547; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  _GEN_780 = 2'h3 == hitsVec_idx ? 1'h0 : _GEN_548; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  _GEN_781 = _sector_hits_T_29 ? _GEN_777 : _GEN_545; // @[TLB.scala 131:34]
  wire  _GEN_782 = _sector_hits_T_29 ? _GEN_778 : _GEN_546; // @[TLB.scala 131:34]
  wire  _GEN_783 = _sector_hits_T_29 ? _GEN_779 : _GEN_547; // @[TLB.scala 131:34]
  wire  _GEN_784 = _sector_hits_T_29 ? _GEN_780 : _GEN_548; // @[TLB.scala 131:34]
  wire  _T_615 = (_sector_hits_T_27[26:18]) == 9'h0; // @[TLB.scala 135:61]
  wire  _GEN_785 = sectored_entries_4_data_0[0] ? 1'h0 : _GEN_781; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  _GEN_786 = sectored_entries_4_data_1[0] ? 1'h0 : _GEN_782; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  _GEN_787 = sectored_entries_4_data_2[0] ? 1'h0 : _GEN_783; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  _GEN_788 = sectored_entries_4_data_3[0] ? 1'h0 : _GEN_784; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  _T_744 = ~(sectored_entries_4_data_0[13]); // @[TLB.scala 143:13]
  wire  _GEN_793 = _T_744 ? 1'h0 : _GEN_545; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _T_745 = ~(sectored_entries_4_data_1[13]); // @[TLB.scala 143:13]
  wire  _GEN_794 = _T_745 ? 1'h0 : _GEN_546; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _T_746 = ~(sectored_entries_4_data_2[13]); // @[TLB.scala 143:13]
  wire  _GEN_795 = _T_746 ? 1'h0 : _GEN_547; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _T_747 = ~(sectored_entries_4_data_3[13]); // @[TLB.scala 143:13]
  wire  _GEN_796 = _T_747 ? 1'h0 : _GEN_548; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _GEN_797 = io_sfence_bits_rs2 & _GEN_793; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _GEN_798 = io_sfence_bits_rs2 & _GEN_794; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _GEN_799 = io_sfence_bits_rs2 & _GEN_795; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _GEN_800 = io_sfence_bits_rs2 & _GEN_796; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _GEN_805 = 2'h0 == hitsVec_idx ? 1'h0 : _GEN_555; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  _GEN_806 = 2'h1 == hitsVec_idx ? 1'h0 : _GEN_556; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  _GEN_807 = 2'h2 == hitsVec_idx ? 1'h0 : _GEN_557; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  _GEN_808 = 2'h3 == hitsVec_idx ? 1'h0 : _GEN_558; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  _GEN_809 = _sector_hits_T_35 ? _GEN_805 : _GEN_555; // @[TLB.scala 131:34]
  wire  _GEN_810 = _sector_hits_T_35 ? _GEN_806 : _GEN_556; // @[TLB.scala 131:34]
  wire  _GEN_811 = _sector_hits_T_35 ? _GEN_807 : _GEN_557; // @[TLB.scala 131:34]
  wire  _GEN_812 = _sector_hits_T_35 ? _GEN_808 : _GEN_558; // @[TLB.scala 131:34]
  wire  _T_754 = (_sector_hits_T_33[26:18]) == 9'h0; // @[TLB.scala 135:61]
  wire  _GEN_813 = sectored_entries_5_data_0[0] ? 1'h0 : _GEN_809; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  _GEN_814 = sectored_entries_5_data_1[0] ? 1'h0 : _GEN_810; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  _GEN_815 = sectored_entries_5_data_2[0] ? 1'h0 : _GEN_811; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  _GEN_816 = sectored_entries_5_data_3[0] ? 1'h0 : _GEN_812; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  _T_883 = ~(sectored_entries_5_data_0[13]); // @[TLB.scala 143:13]
  wire  _GEN_821 = _T_883 ? 1'h0 : _GEN_555; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _T_884 = ~(sectored_entries_5_data_1[13]); // @[TLB.scala 143:13]
  wire  _GEN_822 = _T_884 ? 1'h0 : _GEN_556; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _T_885 = ~(sectored_entries_5_data_2[13]); // @[TLB.scala 143:13]
  wire  _GEN_823 = _T_885 ? 1'h0 : _GEN_557; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _T_886 = ~(sectored_entries_5_data_3[13]); // @[TLB.scala 143:13]
  wire  _GEN_824 = _T_886 ? 1'h0 : _GEN_558; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _GEN_825 = io_sfence_bits_rs2 & _GEN_821; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _GEN_826 = io_sfence_bits_rs2 & _GEN_822; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _GEN_827 = io_sfence_bits_rs2 & _GEN_823; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _GEN_828 = io_sfence_bits_rs2 & _GEN_824; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _GEN_833 = 2'h0 == hitsVec_idx ? 1'h0 : _GEN_565; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  _GEN_834 = 2'h1 == hitsVec_idx ? 1'h0 : _GEN_566; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  _GEN_835 = 2'h2 == hitsVec_idx ? 1'h0 : _GEN_567; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  _GEN_836 = 2'h3 == hitsVec_idx ? 1'h0 : _GEN_568; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  _GEN_837 = _sector_hits_T_41 ? _GEN_833 : _GEN_565; // @[TLB.scala 131:34]
  wire  _GEN_838 = _sector_hits_T_41 ? _GEN_834 : _GEN_566; // @[TLB.scala 131:34]
  wire  _GEN_839 = _sector_hits_T_41 ? _GEN_835 : _GEN_567; // @[TLB.scala 131:34]
  wire  _GEN_840 = _sector_hits_T_41 ? _GEN_836 : _GEN_568; // @[TLB.scala 131:34]
  wire  _T_893 = (_sector_hits_T_39[26:18]) == 9'h0; // @[TLB.scala 135:61]
  wire  _GEN_841 = sectored_entries_6_data_0[0] ? 1'h0 : _GEN_837; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  _GEN_842 = sectored_entries_6_data_1[0] ? 1'h0 : _GEN_838; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  _GEN_843 = sectored_entries_6_data_2[0] ? 1'h0 : _GEN_839; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  _GEN_844 = sectored_entries_6_data_3[0] ? 1'h0 : _GEN_840; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  _T_1022 = ~(sectored_entries_6_data_0[13]); // @[TLB.scala 143:13]
  wire  _GEN_849 = _T_1022 ? 1'h0 : _GEN_565; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _T_1023 = ~(sectored_entries_6_data_1[13]); // @[TLB.scala 143:13]
  wire  _GEN_850 = _T_1023 ? 1'h0 : _GEN_566; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _T_1024 = ~(sectored_entries_6_data_2[13]); // @[TLB.scala 143:13]
  wire  _GEN_851 = _T_1024 ? 1'h0 : _GEN_567; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _T_1025 = ~(sectored_entries_6_data_3[13]); // @[TLB.scala 143:13]
  wire  _GEN_852 = _T_1025 ? 1'h0 : _GEN_568; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _GEN_853 = io_sfence_bits_rs2 & _GEN_849; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _GEN_854 = io_sfence_bits_rs2 & _GEN_850; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _GEN_855 = io_sfence_bits_rs2 & _GEN_851; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _GEN_856 = io_sfence_bits_rs2 & _GEN_852; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _GEN_861 = 2'h0 == hitsVec_idx ? 1'h0 : _GEN_575; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  _GEN_862 = 2'h1 == hitsVec_idx ? 1'h0 : _GEN_576; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  _GEN_863 = 2'h2 == hitsVec_idx ? 1'h0 : _GEN_577; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  _GEN_864 = 2'h3 == hitsVec_idx ? 1'h0 : _GEN_578; // @[TLB.scala 131:58 TLB.scala 131:58]
  wire  _GEN_865 = _sector_hits_T_47 ? _GEN_861 : _GEN_575; // @[TLB.scala 131:34]
  wire  _GEN_866 = _sector_hits_T_47 ? _GEN_862 : _GEN_576; // @[TLB.scala 131:34]
  wire  _GEN_867 = _sector_hits_T_47 ? _GEN_863 : _GEN_577; // @[TLB.scala 131:34]
  wire  _GEN_868 = _sector_hits_T_47 ? _GEN_864 : _GEN_578; // @[TLB.scala 131:34]
  wire  _T_1032 = (_sector_hits_T_45[26:18]) == 9'h0; // @[TLB.scala 135:61]
  wire  _GEN_869 = sectored_entries_7_data_0[0] ? 1'h0 : _GEN_865; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  _GEN_870 = sectored_entries_7_data_1[0] ? 1'h0 : _GEN_866; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  _GEN_871 = sectored_entries_7_data_2[0] ? 1'h0 : _GEN_867; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  _GEN_872 = sectored_entries_7_data_3[0] ? 1'h0 : _GEN_868; // @[TLB.scala 137:41 TLB.scala 137:45]
  wire  _T_1161 = ~(sectored_entries_7_data_0[13]); // @[TLB.scala 143:13]
  wire  _GEN_877 = _T_1161 ? 1'h0 : _GEN_575; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _T_1162 = ~(sectored_entries_7_data_1[13]); // @[TLB.scala 143:13]
  wire  _GEN_878 = _T_1162 ? 1'h0 : _GEN_576; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _T_1163 = ~(sectored_entries_7_data_2[13]); // @[TLB.scala 143:13]
  wire  _GEN_879 = _T_1163 ? 1'h0 : _GEN_577; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _T_1164 = ~(sectored_entries_7_data_3[13]); // @[TLB.scala 143:13]
  wire  _GEN_880 = _T_1164 ? 1'h0 : _GEN_578; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _GEN_881 = io_sfence_bits_rs2 & _GEN_877; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _GEN_882 = io_sfence_bits_rs2 & _GEN_878; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _GEN_883 = io_sfence_bits_rs2 & _GEN_879; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _GEN_884 = io_sfence_bits_rs2 & _GEN_880; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _T_1196 = ~(superpage_entries_0_data_0[13]); // @[TLB.scala 143:13]
  wire  _GEN_890 = _T_1196 ? 1'h0 : _GEN_491; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _GEN_891 = io_sfence_bits_rs2 & _GEN_890; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _T_1228 = ~(superpage_entries_1_data_0[13]); // @[TLB.scala 143:13]
  wire  _GEN_894 = _T_1228 ? 1'h0 : _GEN_495; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _GEN_895 = io_sfence_bits_rs2 & _GEN_894; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _T_1260 = ~(superpage_entries_2_data_0[13]); // @[TLB.scala 143:13]
  wire  _GEN_898 = _T_1260 ? 1'h0 : _GEN_499; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _GEN_899 = io_sfence_bits_rs2 & _GEN_898; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _T_1292 = ~(superpage_entries_3_data_0[13]); // @[TLB.scala 143:13]
  wire  _GEN_902 = _T_1292 ? 1'h0 : _GEN_503; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _GEN_903 = io_sfence_bits_rs2 & _GEN_902; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _T_1324 = ~(special_entry_data_0[13]); // @[TLB.scala 143:13]
  wire  _GEN_906 = _T_1324 ? 1'h0 : _GEN_487; // @[TLB.scala 143:19 TLB.scala 143:23]
  wire  _GEN_907 = io_sfence_bits_rs2 & _GEN_906; // @[TLB.scala 384:40 TLB.scala 126:38]
  wire  _T_1326 = multipleHits | reset; // @[TLB.scala 388:24]
  OptimizationBarrier mpu_ppn_data_barrier ( // @[package.scala 236:25]
    .io_x_ppn(mpu_ppn_data_barrier_io_x_ppn),
    .io_x_u(mpu_ppn_data_barrier_io_x_u),
    .io_x_ae(mpu_ppn_data_barrier_io_x_ae),
    .io_x_sw(mpu_ppn_data_barrier_io_x_sw),
    .io_x_sx(mpu_ppn_data_barrier_io_x_sx),
    .io_x_sr(mpu_ppn_data_barrier_io_x_sr),
    .io_x_pw(mpu_ppn_data_barrier_io_x_pw),
    .io_x_px(mpu_ppn_data_barrier_io_x_px),
    .io_x_pr(mpu_ppn_data_barrier_io_x_pr),
    .io_x_ppp(mpu_ppn_data_barrier_io_x_ppp),
    .io_x_pal(mpu_ppn_data_barrier_io_x_pal),
    .io_x_paa(mpu_ppn_data_barrier_io_x_paa),
    .io_x_eff(mpu_ppn_data_barrier_io_x_eff),
    .io_x_c(mpu_ppn_data_barrier_io_x_c),
    .io_y_ppn(mpu_ppn_data_barrier_io_y_ppn),
    .io_y_u(mpu_ppn_data_barrier_io_y_u),
    .io_y_ae(mpu_ppn_data_barrier_io_y_ae),
    .io_y_sw(mpu_ppn_data_barrier_io_y_sw),
    .io_y_sx(mpu_ppn_data_barrier_io_y_sx),
    .io_y_sr(mpu_ppn_data_barrier_io_y_sr),
    .io_y_pw(mpu_ppn_data_barrier_io_y_pw),
    .io_y_px(mpu_ppn_data_barrier_io_y_px),
    .io_y_pr(mpu_ppn_data_barrier_io_y_pr),
    .io_y_ppp(mpu_ppn_data_barrier_io_y_ppp),
    .io_y_pal(mpu_ppn_data_barrier_io_y_pal),
    .io_y_paa(mpu_ppn_data_barrier_io_y_paa),
    .io_y_eff(mpu_ppn_data_barrier_io_y_eff),
    .io_y_c(mpu_ppn_data_barrier_io_y_c)
  );
  PMPChecker_2 pmp ( // @[TLB.scala 190:19]
    .io_prv(pmp_io_prv),
    .io_pmp_0_cfg_l(pmp_io_pmp_0_cfg_l),
    .io_pmp_0_cfg_a(pmp_io_pmp_0_cfg_a),
    .io_pmp_0_cfg_x(pmp_io_pmp_0_cfg_x),
    .io_pmp_0_cfg_w(pmp_io_pmp_0_cfg_w),
    .io_pmp_0_cfg_r(pmp_io_pmp_0_cfg_r),
    .io_pmp_0_addr(pmp_io_pmp_0_addr),
    .io_pmp_0_mask(pmp_io_pmp_0_mask),
    .io_pmp_1_cfg_l(pmp_io_pmp_1_cfg_l),
    .io_pmp_1_cfg_a(pmp_io_pmp_1_cfg_a),
    .io_pmp_1_cfg_x(pmp_io_pmp_1_cfg_x),
    .io_pmp_1_cfg_w(pmp_io_pmp_1_cfg_w),
    .io_pmp_1_cfg_r(pmp_io_pmp_1_cfg_r),
    .io_pmp_1_addr(pmp_io_pmp_1_addr),
    .io_pmp_1_mask(pmp_io_pmp_1_mask),
    .io_pmp_2_cfg_l(pmp_io_pmp_2_cfg_l),
    .io_pmp_2_cfg_a(pmp_io_pmp_2_cfg_a),
    .io_pmp_2_cfg_x(pmp_io_pmp_2_cfg_x),
    .io_pmp_2_cfg_w(pmp_io_pmp_2_cfg_w),
    .io_pmp_2_cfg_r(pmp_io_pmp_2_cfg_r),
    .io_pmp_2_addr(pmp_io_pmp_2_addr),
    .io_pmp_2_mask(pmp_io_pmp_2_mask),
    .io_pmp_3_cfg_l(pmp_io_pmp_3_cfg_l),
    .io_pmp_3_cfg_a(pmp_io_pmp_3_cfg_a),
    .io_pmp_3_cfg_x(pmp_io_pmp_3_cfg_x),
    .io_pmp_3_cfg_w(pmp_io_pmp_3_cfg_w),
    .io_pmp_3_cfg_r(pmp_io_pmp_3_cfg_r),
    .io_pmp_3_addr(pmp_io_pmp_3_addr),
    .io_pmp_3_mask(pmp_io_pmp_3_mask),
    .io_pmp_4_cfg_l(pmp_io_pmp_4_cfg_l),
    .io_pmp_4_cfg_a(pmp_io_pmp_4_cfg_a),
    .io_pmp_4_cfg_x(pmp_io_pmp_4_cfg_x),
    .io_pmp_4_cfg_w(pmp_io_pmp_4_cfg_w),
    .io_pmp_4_cfg_r(pmp_io_pmp_4_cfg_r),
    .io_pmp_4_addr(pmp_io_pmp_4_addr),
    .io_pmp_4_mask(pmp_io_pmp_4_mask),
    .io_pmp_5_cfg_l(pmp_io_pmp_5_cfg_l),
    .io_pmp_5_cfg_a(pmp_io_pmp_5_cfg_a),
    .io_pmp_5_cfg_x(pmp_io_pmp_5_cfg_x),
    .io_pmp_5_cfg_w(pmp_io_pmp_5_cfg_w),
    .io_pmp_5_cfg_r(pmp_io_pmp_5_cfg_r),
    .io_pmp_5_addr(pmp_io_pmp_5_addr),
    .io_pmp_5_mask(pmp_io_pmp_5_mask),
    .io_pmp_6_cfg_l(pmp_io_pmp_6_cfg_l),
    .io_pmp_6_cfg_a(pmp_io_pmp_6_cfg_a),
    .io_pmp_6_cfg_x(pmp_io_pmp_6_cfg_x),
    .io_pmp_6_cfg_w(pmp_io_pmp_6_cfg_w),
    .io_pmp_6_cfg_r(pmp_io_pmp_6_cfg_r),
    .io_pmp_6_addr(pmp_io_pmp_6_addr),
    .io_pmp_6_mask(pmp_io_pmp_6_mask),
    .io_pmp_7_cfg_l(pmp_io_pmp_7_cfg_l),
    .io_pmp_7_cfg_a(pmp_io_pmp_7_cfg_a),
    .io_pmp_7_cfg_x(pmp_io_pmp_7_cfg_x),
    .io_pmp_7_cfg_w(pmp_io_pmp_7_cfg_w),
    .io_pmp_7_cfg_r(pmp_io_pmp_7_cfg_r),
    .io_pmp_7_addr(pmp_io_pmp_7_addr),
    .io_pmp_7_mask(pmp_io_pmp_7_mask),
    .io_addr(pmp_io_addr),
    .io_r(pmp_io_r),
    .io_w(pmp_io_w),
    .io_x(pmp_io_x)
  );
  OptimizationBarrier ppn_data_barrier ( // @[package.scala 236:25]
    .io_x_ppn(ppn_data_barrier_io_x_ppn),
    .io_x_u(ppn_data_barrier_io_x_u),
    .io_x_ae(ppn_data_barrier_io_x_ae),
    .io_x_sw(ppn_data_barrier_io_x_sw),
    .io_x_sx(ppn_data_barrier_io_x_sx),
    .io_x_sr(ppn_data_barrier_io_x_sr),
    .io_x_pw(ppn_data_barrier_io_x_pw),
    .io_x_px(ppn_data_barrier_io_x_px),
    .io_x_pr(ppn_data_barrier_io_x_pr),
    .io_x_ppp(ppn_data_barrier_io_x_ppp),
    .io_x_pal(ppn_data_barrier_io_x_pal),
    .io_x_paa(ppn_data_barrier_io_x_paa),
    .io_x_eff(ppn_data_barrier_io_x_eff),
    .io_x_c(ppn_data_barrier_io_x_c),
    .io_y_ppn(ppn_data_barrier_io_y_ppn),
    .io_y_u(ppn_data_barrier_io_y_u),
    .io_y_ae(ppn_data_barrier_io_y_ae),
    .io_y_sw(ppn_data_barrier_io_y_sw),
    .io_y_sx(ppn_data_barrier_io_y_sx),
    .io_y_sr(ppn_data_barrier_io_y_sr),
    .io_y_pw(ppn_data_barrier_io_y_pw),
    .io_y_px(ppn_data_barrier_io_y_px),
    .io_y_pr(ppn_data_barrier_io_y_pr),
    .io_y_ppp(ppn_data_barrier_io_y_ppp),
    .io_y_pal(ppn_data_barrier_io_y_pal),
    .io_y_paa(ppn_data_barrier_io_y_paa),
    .io_y_eff(ppn_data_barrier_io_y_eff),
    .io_y_c(ppn_data_barrier_io_y_c)
  );
  OptimizationBarrier ppn_data_barrier_1 ( // @[package.scala 236:25]
    .io_x_ppn(ppn_data_barrier_1_io_x_ppn),
    .io_x_u(ppn_data_barrier_1_io_x_u),
    .io_x_ae(ppn_data_barrier_1_io_x_ae),
    .io_x_sw(ppn_data_barrier_1_io_x_sw),
    .io_x_sx(ppn_data_barrier_1_io_x_sx),
    .io_x_sr(ppn_data_barrier_1_io_x_sr),
    .io_x_pw(ppn_data_barrier_1_io_x_pw),
    .io_x_px(ppn_data_barrier_1_io_x_px),
    .io_x_pr(ppn_data_barrier_1_io_x_pr),
    .io_x_ppp(ppn_data_barrier_1_io_x_ppp),
    .io_x_pal(ppn_data_barrier_1_io_x_pal),
    .io_x_paa(ppn_data_barrier_1_io_x_paa),
    .io_x_eff(ppn_data_barrier_1_io_x_eff),
    .io_x_c(ppn_data_barrier_1_io_x_c),
    .io_y_ppn(ppn_data_barrier_1_io_y_ppn),
    .io_y_u(ppn_data_barrier_1_io_y_u),
    .io_y_ae(ppn_data_barrier_1_io_y_ae),
    .io_y_sw(ppn_data_barrier_1_io_y_sw),
    .io_y_sx(ppn_data_barrier_1_io_y_sx),
    .io_y_sr(ppn_data_barrier_1_io_y_sr),
    .io_y_pw(ppn_data_barrier_1_io_y_pw),
    .io_y_px(ppn_data_barrier_1_io_y_px),
    .io_y_pr(ppn_data_barrier_1_io_y_pr),
    .io_y_ppp(ppn_data_barrier_1_io_y_ppp),
    .io_y_pal(ppn_data_barrier_1_io_y_pal),
    .io_y_paa(ppn_data_barrier_1_io_y_paa),
    .io_y_eff(ppn_data_barrier_1_io_y_eff),
    .io_y_c(ppn_data_barrier_1_io_y_c)
  );
  OptimizationBarrier ppn_data_barrier_2 ( // @[package.scala 236:25]
    .io_x_ppn(ppn_data_barrier_2_io_x_ppn),
    .io_x_u(ppn_data_barrier_2_io_x_u),
    .io_x_ae(ppn_data_barrier_2_io_x_ae),
    .io_x_sw(ppn_data_barrier_2_io_x_sw),
    .io_x_sx(ppn_data_barrier_2_io_x_sx),
    .io_x_sr(ppn_data_barrier_2_io_x_sr),
    .io_x_pw(ppn_data_barrier_2_io_x_pw),
    .io_x_px(ppn_data_barrier_2_io_x_px),
    .io_x_pr(ppn_data_barrier_2_io_x_pr),
    .io_x_ppp(ppn_data_barrier_2_io_x_ppp),
    .io_x_pal(ppn_data_barrier_2_io_x_pal),
    .io_x_paa(ppn_data_barrier_2_io_x_paa),
    .io_x_eff(ppn_data_barrier_2_io_x_eff),
    .io_x_c(ppn_data_barrier_2_io_x_c),
    .io_y_ppn(ppn_data_barrier_2_io_y_ppn),
    .io_y_u(ppn_data_barrier_2_io_y_u),
    .io_y_ae(ppn_data_barrier_2_io_y_ae),
    .io_y_sw(ppn_data_barrier_2_io_y_sw),
    .io_y_sx(ppn_data_barrier_2_io_y_sx),
    .io_y_sr(ppn_data_barrier_2_io_y_sr),
    .io_y_pw(ppn_data_barrier_2_io_y_pw),
    .io_y_px(ppn_data_barrier_2_io_y_px),
    .io_y_pr(ppn_data_barrier_2_io_y_pr),
    .io_y_ppp(ppn_data_barrier_2_io_y_ppp),
    .io_y_pal(ppn_data_barrier_2_io_y_pal),
    .io_y_paa(ppn_data_barrier_2_io_y_paa),
    .io_y_eff(ppn_data_barrier_2_io_y_eff),
    .io_y_c(ppn_data_barrier_2_io_y_c)
  );
  OptimizationBarrier ppn_data_barrier_3 ( // @[package.scala 236:25]
    .io_x_ppn(ppn_data_barrier_3_io_x_ppn),
    .io_x_u(ppn_data_barrier_3_io_x_u),
    .io_x_ae(ppn_data_barrier_3_io_x_ae),
    .io_x_sw(ppn_data_barrier_3_io_x_sw),
    .io_x_sx(ppn_data_barrier_3_io_x_sx),
    .io_x_sr(ppn_data_barrier_3_io_x_sr),
    .io_x_pw(ppn_data_barrier_3_io_x_pw),
    .io_x_px(ppn_data_barrier_3_io_x_px),
    .io_x_pr(ppn_data_barrier_3_io_x_pr),
    .io_x_ppp(ppn_data_barrier_3_io_x_ppp),
    .io_x_pal(ppn_data_barrier_3_io_x_pal),
    .io_x_paa(ppn_data_barrier_3_io_x_paa),
    .io_x_eff(ppn_data_barrier_3_io_x_eff),
    .io_x_c(ppn_data_barrier_3_io_x_c),
    .io_y_ppn(ppn_data_barrier_3_io_y_ppn),
    .io_y_u(ppn_data_barrier_3_io_y_u),
    .io_y_ae(ppn_data_barrier_3_io_y_ae),
    .io_y_sw(ppn_data_barrier_3_io_y_sw),
    .io_y_sx(ppn_data_barrier_3_io_y_sx),
    .io_y_sr(ppn_data_barrier_3_io_y_sr),
    .io_y_pw(ppn_data_barrier_3_io_y_pw),
    .io_y_px(ppn_data_barrier_3_io_y_px),
    .io_y_pr(ppn_data_barrier_3_io_y_pr),
    .io_y_ppp(ppn_data_barrier_3_io_y_ppp),
    .io_y_pal(ppn_data_barrier_3_io_y_pal),
    .io_y_paa(ppn_data_barrier_3_io_y_paa),
    .io_y_eff(ppn_data_barrier_3_io_y_eff),
    .io_y_c(ppn_data_barrier_3_io_y_c)
  );
  OptimizationBarrier ppn_data_barrier_4 ( // @[package.scala 236:25]
    .io_x_ppn(ppn_data_barrier_4_io_x_ppn),
    .io_x_u(ppn_data_barrier_4_io_x_u),
    .io_x_ae(ppn_data_barrier_4_io_x_ae),
    .io_x_sw(ppn_data_barrier_4_io_x_sw),
    .io_x_sx(ppn_data_barrier_4_io_x_sx),
    .io_x_sr(ppn_data_barrier_4_io_x_sr),
    .io_x_pw(ppn_data_barrier_4_io_x_pw),
    .io_x_px(ppn_data_barrier_4_io_x_px),
    .io_x_pr(ppn_data_barrier_4_io_x_pr),
    .io_x_ppp(ppn_data_barrier_4_io_x_ppp),
    .io_x_pal(ppn_data_barrier_4_io_x_pal),
    .io_x_paa(ppn_data_barrier_4_io_x_paa),
    .io_x_eff(ppn_data_barrier_4_io_x_eff),
    .io_x_c(ppn_data_barrier_4_io_x_c),
    .io_y_ppn(ppn_data_barrier_4_io_y_ppn),
    .io_y_u(ppn_data_barrier_4_io_y_u),
    .io_y_ae(ppn_data_barrier_4_io_y_ae),
    .io_y_sw(ppn_data_barrier_4_io_y_sw),
    .io_y_sx(ppn_data_barrier_4_io_y_sx),
    .io_y_sr(ppn_data_barrier_4_io_y_sr),
    .io_y_pw(ppn_data_barrier_4_io_y_pw),
    .io_y_px(ppn_data_barrier_4_io_y_px),
    .io_y_pr(ppn_data_barrier_4_io_y_pr),
    .io_y_ppp(ppn_data_barrier_4_io_y_ppp),
    .io_y_pal(ppn_data_barrier_4_io_y_pal),
    .io_y_paa(ppn_data_barrier_4_io_y_paa),
    .io_y_eff(ppn_data_barrier_4_io_y_eff),
    .io_y_c(ppn_data_barrier_4_io_y_c)
  );
  OptimizationBarrier ppn_data_barrier_5 ( // @[package.scala 236:25]
    .io_x_ppn(ppn_data_barrier_5_io_x_ppn),
    .io_x_u(ppn_data_barrier_5_io_x_u),
    .io_x_ae(ppn_data_barrier_5_io_x_ae),
    .io_x_sw(ppn_data_barrier_5_io_x_sw),
    .io_x_sx(ppn_data_barrier_5_io_x_sx),
    .io_x_sr(ppn_data_barrier_5_io_x_sr),
    .io_x_pw(ppn_data_barrier_5_io_x_pw),
    .io_x_px(ppn_data_barrier_5_io_x_px),
    .io_x_pr(ppn_data_barrier_5_io_x_pr),
    .io_x_ppp(ppn_data_barrier_5_io_x_ppp),
    .io_x_pal(ppn_data_barrier_5_io_x_pal),
    .io_x_paa(ppn_data_barrier_5_io_x_paa),
    .io_x_eff(ppn_data_barrier_5_io_x_eff),
    .io_x_c(ppn_data_barrier_5_io_x_c),
    .io_y_ppn(ppn_data_barrier_5_io_y_ppn),
    .io_y_u(ppn_data_barrier_5_io_y_u),
    .io_y_ae(ppn_data_barrier_5_io_y_ae),
    .io_y_sw(ppn_data_barrier_5_io_y_sw),
    .io_y_sx(ppn_data_barrier_5_io_y_sx),
    .io_y_sr(ppn_data_barrier_5_io_y_sr),
    .io_y_pw(ppn_data_barrier_5_io_y_pw),
    .io_y_px(ppn_data_barrier_5_io_y_px),
    .io_y_pr(ppn_data_barrier_5_io_y_pr),
    .io_y_ppp(ppn_data_barrier_5_io_y_ppp),
    .io_y_pal(ppn_data_barrier_5_io_y_pal),
    .io_y_paa(ppn_data_barrier_5_io_y_paa),
    .io_y_eff(ppn_data_barrier_5_io_y_eff),
    .io_y_c(ppn_data_barrier_5_io_y_c)
  );
  OptimizationBarrier ppn_data_barrier_6 ( // @[package.scala 236:25]
    .io_x_ppn(ppn_data_barrier_6_io_x_ppn),
    .io_x_u(ppn_data_barrier_6_io_x_u),
    .io_x_ae(ppn_data_barrier_6_io_x_ae),
    .io_x_sw(ppn_data_barrier_6_io_x_sw),
    .io_x_sx(ppn_data_barrier_6_io_x_sx),
    .io_x_sr(ppn_data_barrier_6_io_x_sr),
    .io_x_pw(ppn_data_barrier_6_io_x_pw),
    .io_x_px(ppn_data_barrier_6_io_x_px),
    .io_x_pr(ppn_data_barrier_6_io_x_pr),
    .io_x_ppp(ppn_data_barrier_6_io_x_ppp),
    .io_x_pal(ppn_data_barrier_6_io_x_pal),
    .io_x_paa(ppn_data_barrier_6_io_x_paa),
    .io_x_eff(ppn_data_barrier_6_io_x_eff),
    .io_x_c(ppn_data_barrier_6_io_x_c),
    .io_y_ppn(ppn_data_barrier_6_io_y_ppn),
    .io_y_u(ppn_data_barrier_6_io_y_u),
    .io_y_ae(ppn_data_barrier_6_io_y_ae),
    .io_y_sw(ppn_data_barrier_6_io_y_sw),
    .io_y_sx(ppn_data_barrier_6_io_y_sx),
    .io_y_sr(ppn_data_barrier_6_io_y_sr),
    .io_y_pw(ppn_data_barrier_6_io_y_pw),
    .io_y_px(ppn_data_barrier_6_io_y_px),
    .io_y_pr(ppn_data_barrier_6_io_y_pr),
    .io_y_ppp(ppn_data_barrier_6_io_y_ppp),
    .io_y_pal(ppn_data_barrier_6_io_y_pal),
    .io_y_paa(ppn_data_barrier_6_io_y_paa),
    .io_y_eff(ppn_data_barrier_6_io_y_eff),
    .io_y_c(ppn_data_barrier_6_io_y_c)
  );
  OptimizationBarrier ppn_data_barrier_7 ( // @[package.scala 236:25]
    .io_x_ppn(ppn_data_barrier_7_io_x_ppn),
    .io_x_u(ppn_data_barrier_7_io_x_u),
    .io_x_ae(ppn_data_barrier_7_io_x_ae),
    .io_x_sw(ppn_data_barrier_7_io_x_sw),
    .io_x_sx(ppn_data_barrier_7_io_x_sx),
    .io_x_sr(ppn_data_barrier_7_io_x_sr),
    .io_x_pw(ppn_data_barrier_7_io_x_pw),
    .io_x_px(ppn_data_barrier_7_io_x_px),
    .io_x_pr(ppn_data_barrier_7_io_x_pr),
    .io_x_ppp(ppn_data_barrier_7_io_x_ppp),
    .io_x_pal(ppn_data_barrier_7_io_x_pal),
    .io_x_paa(ppn_data_barrier_7_io_x_paa),
    .io_x_eff(ppn_data_barrier_7_io_x_eff),
    .io_x_c(ppn_data_barrier_7_io_x_c),
    .io_y_ppn(ppn_data_barrier_7_io_y_ppn),
    .io_y_u(ppn_data_barrier_7_io_y_u),
    .io_y_ae(ppn_data_barrier_7_io_y_ae),
    .io_y_sw(ppn_data_barrier_7_io_y_sw),
    .io_y_sx(ppn_data_barrier_7_io_y_sx),
    .io_y_sr(ppn_data_barrier_7_io_y_sr),
    .io_y_pw(ppn_data_barrier_7_io_y_pw),
    .io_y_px(ppn_data_barrier_7_io_y_px),
    .io_y_pr(ppn_data_barrier_7_io_y_pr),
    .io_y_ppp(ppn_data_barrier_7_io_y_ppp),
    .io_y_pal(ppn_data_barrier_7_io_y_pal),
    .io_y_paa(ppn_data_barrier_7_io_y_paa),
    .io_y_eff(ppn_data_barrier_7_io_y_eff),
    .io_y_c(ppn_data_barrier_7_io_y_c)
  );
  OptimizationBarrier ppn_data_barrier_8 ( // @[package.scala 236:25]
    .io_x_ppn(ppn_data_barrier_8_io_x_ppn),
    .io_x_u(ppn_data_barrier_8_io_x_u),
    .io_x_ae(ppn_data_barrier_8_io_x_ae),
    .io_x_sw(ppn_data_barrier_8_io_x_sw),
    .io_x_sx(ppn_data_barrier_8_io_x_sx),
    .io_x_sr(ppn_data_barrier_8_io_x_sr),
    .io_x_pw(ppn_data_barrier_8_io_x_pw),
    .io_x_px(ppn_data_barrier_8_io_x_px),
    .io_x_pr(ppn_data_barrier_8_io_x_pr),
    .io_x_ppp(ppn_data_barrier_8_io_x_ppp),
    .io_x_pal(ppn_data_barrier_8_io_x_pal),
    .io_x_paa(ppn_data_barrier_8_io_x_paa),
    .io_x_eff(ppn_data_barrier_8_io_x_eff),
    .io_x_c(ppn_data_barrier_8_io_x_c),
    .io_y_ppn(ppn_data_barrier_8_io_y_ppn),
    .io_y_u(ppn_data_barrier_8_io_y_u),
    .io_y_ae(ppn_data_barrier_8_io_y_ae),
    .io_y_sw(ppn_data_barrier_8_io_y_sw),
    .io_y_sx(ppn_data_barrier_8_io_y_sx),
    .io_y_sr(ppn_data_barrier_8_io_y_sr),
    .io_y_pw(ppn_data_barrier_8_io_y_pw),
    .io_y_px(ppn_data_barrier_8_io_y_px),
    .io_y_pr(ppn_data_barrier_8_io_y_pr),
    .io_y_ppp(ppn_data_barrier_8_io_y_ppp),
    .io_y_pal(ppn_data_barrier_8_io_y_pal),
    .io_y_paa(ppn_data_barrier_8_io_y_paa),
    .io_y_eff(ppn_data_barrier_8_io_y_eff),
    .io_y_c(ppn_data_barrier_8_io_y_c)
  );
  OptimizationBarrier ppn_data_barrier_9 ( // @[package.scala 236:25]
    .io_x_ppn(ppn_data_barrier_9_io_x_ppn),
    .io_x_u(ppn_data_barrier_9_io_x_u),
    .io_x_ae(ppn_data_barrier_9_io_x_ae),
    .io_x_sw(ppn_data_barrier_9_io_x_sw),
    .io_x_sx(ppn_data_barrier_9_io_x_sx),
    .io_x_sr(ppn_data_barrier_9_io_x_sr),
    .io_x_pw(ppn_data_barrier_9_io_x_pw),
    .io_x_px(ppn_data_barrier_9_io_x_px),
    .io_x_pr(ppn_data_barrier_9_io_x_pr),
    .io_x_ppp(ppn_data_barrier_9_io_x_ppp),
    .io_x_pal(ppn_data_barrier_9_io_x_pal),
    .io_x_paa(ppn_data_barrier_9_io_x_paa),
    .io_x_eff(ppn_data_barrier_9_io_x_eff),
    .io_x_c(ppn_data_barrier_9_io_x_c),
    .io_y_ppn(ppn_data_barrier_9_io_y_ppn),
    .io_y_u(ppn_data_barrier_9_io_y_u),
    .io_y_ae(ppn_data_barrier_9_io_y_ae),
    .io_y_sw(ppn_data_barrier_9_io_y_sw),
    .io_y_sx(ppn_data_barrier_9_io_y_sx),
    .io_y_sr(ppn_data_barrier_9_io_y_sr),
    .io_y_pw(ppn_data_barrier_9_io_y_pw),
    .io_y_px(ppn_data_barrier_9_io_y_px),
    .io_y_pr(ppn_data_barrier_9_io_y_pr),
    .io_y_ppp(ppn_data_barrier_9_io_y_ppp),
    .io_y_pal(ppn_data_barrier_9_io_y_pal),
    .io_y_paa(ppn_data_barrier_9_io_y_paa),
    .io_y_eff(ppn_data_barrier_9_io_y_eff),
    .io_y_c(ppn_data_barrier_9_io_y_c)
  );
  OptimizationBarrier ppn_data_barrier_10 ( // @[package.scala 236:25]
    .io_x_ppn(ppn_data_barrier_10_io_x_ppn),
    .io_x_u(ppn_data_barrier_10_io_x_u),
    .io_x_ae(ppn_data_barrier_10_io_x_ae),
    .io_x_sw(ppn_data_barrier_10_io_x_sw),
    .io_x_sx(ppn_data_barrier_10_io_x_sx),
    .io_x_sr(ppn_data_barrier_10_io_x_sr),
    .io_x_pw(ppn_data_barrier_10_io_x_pw),
    .io_x_px(ppn_data_barrier_10_io_x_px),
    .io_x_pr(ppn_data_barrier_10_io_x_pr),
    .io_x_ppp(ppn_data_barrier_10_io_x_ppp),
    .io_x_pal(ppn_data_barrier_10_io_x_pal),
    .io_x_paa(ppn_data_barrier_10_io_x_paa),
    .io_x_eff(ppn_data_barrier_10_io_x_eff),
    .io_x_c(ppn_data_barrier_10_io_x_c),
    .io_y_ppn(ppn_data_barrier_10_io_y_ppn),
    .io_y_u(ppn_data_barrier_10_io_y_u),
    .io_y_ae(ppn_data_barrier_10_io_y_ae),
    .io_y_sw(ppn_data_barrier_10_io_y_sw),
    .io_y_sx(ppn_data_barrier_10_io_y_sx),
    .io_y_sr(ppn_data_barrier_10_io_y_sr),
    .io_y_pw(ppn_data_barrier_10_io_y_pw),
    .io_y_px(ppn_data_barrier_10_io_y_px),
    .io_y_pr(ppn_data_barrier_10_io_y_pr),
    .io_y_ppp(ppn_data_barrier_10_io_y_ppp),
    .io_y_pal(ppn_data_barrier_10_io_y_pal),
    .io_y_paa(ppn_data_barrier_10_io_y_paa),
    .io_y_eff(ppn_data_barrier_10_io_y_eff),
    .io_y_c(ppn_data_barrier_10_io_y_c)
  );
  OptimizationBarrier ppn_data_barrier_11 ( // @[package.scala 236:25]
    .io_x_ppn(ppn_data_barrier_11_io_x_ppn),
    .io_x_u(ppn_data_barrier_11_io_x_u),
    .io_x_ae(ppn_data_barrier_11_io_x_ae),
    .io_x_sw(ppn_data_barrier_11_io_x_sw),
    .io_x_sx(ppn_data_barrier_11_io_x_sx),
    .io_x_sr(ppn_data_barrier_11_io_x_sr),
    .io_x_pw(ppn_data_barrier_11_io_x_pw),
    .io_x_px(ppn_data_barrier_11_io_x_px),
    .io_x_pr(ppn_data_barrier_11_io_x_pr),
    .io_x_ppp(ppn_data_barrier_11_io_x_ppp),
    .io_x_pal(ppn_data_barrier_11_io_x_pal),
    .io_x_paa(ppn_data_barrier_11_io_x_paa),
    .io_x_eff(ppn_data_barrier_11_io_x_eff),
    .io_x_c(ppn_data_barrier_11_io_x_c),
    .io_y_ppn(ppn_data_barrier_11_io_y_ppn),
    .io_y_u(ppn_data_barrier_11_io_y_u),
    .io_y_ae(ppn_data_barrier_11_io_y_ae),
    .io_y_sw(ppn_data_barrier_11_io_y_sw),
    .io_y_sx(ppn_data_barrier_11_io_y_sx),
    .io_y_sr(ppn_data_barrier_11_io_y_sr),
    .io_y_pw(ppn_data_barrier_11_io_y_pw),
    .io_y_px(ppn_data_barrier_11_io_y_px),
    .io_y_pr(ppn_data_barrier_11_io_y_pr),
    .io_y_ppp(ppn_data_barrier_11_io_y_ppp),
    .io_y_pal(ppn_data_barrier_11_io_y_pal),
    .io_y_paa(ppn_data_barrier_11_io_y_paa),
    .io_y_eff(ppn_data_barrier_11_io_y_eff),
    .io_y_c(ppn_data_barrier_11_io_y_c)
  );
  OptimizationBarrier ppn_data_barrier_12 ( // @[package.scala 236:25]
    .io_x_ppn(ppn_data_barrier_12_io_x_ppn),
    .io_x_u(ppn_data_barrier_12_io_x_u),
    .io_x_ae(ppn_data_barrier_12_io_x_ae),
    .io_x_sw(ppn_data_barrier_12_io_x_sw),
    .io_x_sx(ppn_data_barrier_12_io_x_sx),
    .io_x_sr(ppn_data_barrier_12_io_x_sr),
    .io_x_pw(ppn_data_barrier_12_io_x_pw),
    .io_x_px(ppn_data_barrier_12_io_x_px),
    .io_x_pr(ppn_data_barrier_12_io_x_pr),
    .io_x_ppp(ppn_data_barrier_12_io_x_ppp),
    .io_x_pal(ppn_data_barrier_12_io_x_pal),
    .io_x_paa(ppn_data_barrier_12_io_x_paa),
    .io_x_eff(ppn_data_barrier_12_io_x_eff),
    .io_x_c(ppn_data_barrier_12_io_x_c),
    .io_y_ppn(ppn_data_barrier_12_io_y_ppn),
    .io_y_u(ppn_data_barrier_12_io_y_u),
    .io_y_ae(ppn_data_barrier_12_io_y_ae),
    .io_y_sw(ppn_data_barrier_12_io_y_sw),
    .io_y_sx(ppn_data_barrier_12_io_y_sx),
    .io_y_sr(ppn_data_barrier_12_io_y_sr),
    .io_y_pw(ppn_data_barrier_12_io_y_pw),
    .io_y_px(ppn_data_barrier_12_io_y_px),
    .io_y_pr(ppn_data_barrier_12_io_y_pr),
    .io_y_ppp(ppn_data_barrier_12_io_y_ppp),
    .io_y_pal(ppn_data_barrier_12_io_y_pal),
    .io_y_paa(ppn_data_barrier_12_io_y_paa),
    .io_y_eff(ppn_data_barrier_12_io_y_eff),
    .io_y_c(ppn_data_barrier_12_io_y_c)
  );
  OptimizationBarrier entries_barrier ( // @[package.scala 236:25]
    .io_x_ppn(entries_barrier_io_x_ppn),
    .io_x_u(entries_barrier_io_x_u),
    .io_x_ae(entries_barrier_io_x_ae),
    .io_x_sw(entries_barrier_io_x_sw),
    .io_x_sx(entries_barrier_io_x_sx),
    .io_x_sr(entries_barrier_io_x_sr),
    .io_x_pw(entries_barrier_io_x_pw),
    .io_x_px(entries_barrier_io_x_px),
    .io_x_pr(entries_barrier_io_x_pr),
    .io_x_ppp(entries_barrier_io_x_ppp),
    .io_x_pal(entries_barrier_io_x_pal),
    .io_x_paa(entries_barrier_io_x_paa),
    .io_x_eff(entries_barrier_io_x_eff),
    .io_x_c(entries_barrier_io_x_c),
    .io_y_ppn(entries_barrier_io_y_ppn),
    .io_y_u(entries_barrier_io_y_u),
    .io_y_ae(entries_barrier_io_y_ae),
    .io_y_sw(entries_barrier_io_y_sw),
    .io_y_sx(entries_barrier_io_y_sx),
    .io_y_sr(entries_barrier_io_y_sr),
    .io_y_pw(entries_barrier_io_y_pw),
    .io_y_px(entries_barrier_io_y_px),
    .io_y_pr(entries_barrier_io_y_pr),
    .io_y_ppp(entries_barrier_io_y_ppp),
    .io_y_pal(entries_barrier_io_y_pal),
    .io_y_paa(entries_barrier_io_y_paa),
    .io_y_eff(entries_barrier_io_y_eff),
    .io_y_c(entries_barrier_io_y_c)
  );
  OptimizationBarrier entries_barrier_1 ( // @[package.scala 236:25]
    .io_x_ppn(entries_barrier_1_io_x_ppn),
    .io_x_u(entries_barrier_1_io_x_u),
    .io_x_ae(entries_barrier_1_io_x_ae),
    .io_x_sw(entries_barrier_1_io_x_sw),
    .io_x_sx(entries_barrier_1_io_x_sx),
    .io_x_sr(entries_barrier_1_io_x_sr),
    .io_x_pw(entries_barrier_1_io_x_pw),
    .io_x_px(entries_barrier_1_io_x_px),
    .io_x_pr(entries_barrier_1_io_x_pr),
    .io_x_ppp(entries_barrier_1_io_x_ppp),
    .io_x_pal(entries_barrier_1_io_x_pal),
    .io_x_paa(entries_barrier_1_io_x_paa),
    .io_x_eff(entries_barrier_1_io_x_eff),
    .io_x_c(entries_barrier_1_io_x_c),
    .io_y_ppn(entries_barrier_1_io_y_ppn),
    .io_y_u(entries_barrier_1_io_y_u),
    .io_y_ae(entries_barrier_1_io_y_ae),
    .io_y_sw(entries_barrier_1_io_y_sw),
    .io_y_sx(entries_barrier_1_io_y_sx),
    .io_y_sr(entries_barrier_1_io_y_sr),
    .io_y_pw(entries_barrier_1_io_y_pw),
    .io_y_px(entries_barrier_1_io_y_px),
    .io_y_pr(entries_barrier_1_io_y_pr),
    .io_y_ppp(entries_barrier_1_io_y_ppp),
    .io_y_pal(entries_barrier_1_io_y_pal),
    .io_y_paa(entries_barrier_1_io_y_paa),
    .io_y_eff(entries_barrier_1_io_y_eff),
    .io_y_c(entries_barrier_1_io_y_c)
  );
  OptimizationBarrier entries_barrier_2 ( // @[package.scala 236:25]
    .io_x_ppn(entries_barrier_2_io_x_ppn),
    .io_x_u(entries_barrier_2_io_x_u),
    .io_x_ae(entries_barrier_2_io_x_ae),
    .io_x_sw(entries_barrier_2_io_x_sw),
    .io_x_sx(entries_barrier_2_io_x_sx),
    .io_x_sr(entries_barrier_2_io_x_sr),
    .io_x_pw(entries_barrier_2_io_x_pw),
    .io_x_px(entries_barrier_2_io_x_px),
    .io_x_pr(entries_barrier_2_io_x_pr),
    .io_x_ppp(entries_barrier_2_io_x_ppp),
    .io_x_pal(entries_barrier_2_io_x_pal),
    .io_x_paa(entries_barrier_2_io_x_paa),
    .io_x_eff(entries_barrier_2_io_x_eff),
    .io_x_c(entries_barrier_2_io_x_c),
    .io_y_ppn(entries_barrier_2_io_y_ppn),
    .io_y_u(entries_barrier_2_io_y_u),
    .io_y_ae(entries_barrier_2_io_y_ae),
    .io_y_sw(entries_barrier_2_io_y_sw),
    .io_y_sx(entries_barrier_2_io_y_sx),
    .io_y_sr(entries_barrier_2_io_y_sr),
    .io_y_pw(entries_barrier_2_io_y_pw),
    .io_y_px(entries_barrier_2_io_y_px),
    .io_y_pr(entries_barrier_2_io_y_pr),
    .io_y_ppp(entries_barrier_2_io_y_ppp),
    .io_y_pal(entries_barrier_2_io_y_pal),
    .io_y_paa(entries_barrier_2_io_y_paa),
    .io_y_eff(entries_barrier_2_io_y_eff),
    .io_y_c(entries_barrier_2_io_y_c)
  );
  OptimizationBarrier entries_barrier_3 ( // @[package.scala 236:25]
    .io_x_ppn(entries_barrier_3_io_x_ppn),
    .io_x_u(entries_barrier_3_io_x_u),
    .io_x_ae(entries_barrier_3_io_x_ae),
    .io_x_sw(entries_barrier_3_io_x_sw),
    .io_x_sx(entries_barrier_3_io_x_sx),
    .io_x_sr(entries_barrier_3_io_x_sr),
    .io_x_pw(entries_barrier_3_io_x_pw),
    .io_x_px(entries_barrier_3_io_x_px),
    .io_x_pr(entries_barrier_3_io_x_pr),
    .io_x_ppp(entries_barrier_3_io_x_ppp),
    .io_x_pal(entries_barrier_3_io_x_pal),
    .io_x_paa(entries_barrier_3_io_x_paa),
    .io_x_eff(entries_barrier_3_io_x_eff),
    .io_x_c(entries_barrier_3_io_x_c),
    .io_y_ppn(entries_barrier_3_io_y_ppn),
    .io_y_u(entries_barrier_3_io_y_u),
    .io_y_ae(entries_barrier_3_io_y_ae),
    .io_y_sw(entries_barrier_3_io_y_sw),
    .io_y_sx(entries_barrier_3_io_y_sx),
    .io_y_sr(entries_barrier_3_io_y_sr),
    .io_y_pw(entries_barrier_3_io_y_pw),
    .io_y_px(entries_barrier_3_io_y_px),
    .io_y_pr(entries_barrier_3_io_y_pr),
    .io_y_ppp(entries_barrier_3_io_y_ppp),
    .io_y_pal(entries_barrier_3_io_y_pal),
    .io_y_paa(entries_barrier_3_io_y_paa),
    .io_y_eff(entries_barrier_3_io_y_eff),
    .io_y_c(entries_barrier_3_io_y_c)
  );
  OptimizationBarrier entries_barrier_4 ( // @[package.scala 236:25]
    .io_x_ppn(entries_barrier_4_io_x_ppn),
    .io_x_u(entries_barrier_4_io_x_u),
    .io_x_ae(entries_barrier_4_io_x_ae),
    .io_x_sw(entries_barrier_4_io_x_sw),
    .io_x_sx(entries_barrier_4_io_x_sx),
    .io_x_sr(entries_barrier_4_io_x_sr),
    .io_x_pw(entries_barrier_4_io_x_pw),
    .io_x_px(entries_barrier_4_io_x_px),
    .io_x_pr(entries_barrier_4_io_x_pr),
    .io_x_ppp(entries_barrier_4_io_x_ppp),
    .io_x_pal(entries_barrier_4_io_x_pal),
    .io_x_paa(entries_barrier_4_io_x_paa),
    .io_x_eff(entries_barrier_4_io_x_eff),
    .io_x_c(entries_barrier_4_io_x_c),
    .io_y_ppn(entries_barrier_4_io_y_ppn),
    .io_y_u(entries_barrier_4_io_y_u),
    .io_y_ae(entries_barrier_4_io_y_ae),
    .io_y_sw(entries_barrier_4_io_y_sw),
    .io_y_sx(entries_barrier_4_io_y_sx),
    .io_y_sr(entries_barrier_4_io_y_sr),
    .io_y_pw(entries_barrier_4_io_y_pw),
    .io_y_px(entries_barrier_4_io_y_px),
    .io_y_pr(entries_barrier_4_io_y_pr),
    .io_y_ppp(entries_barrier_4_io_y_ppp),
    .io_y_pal(entries_barrier_4_io_y_pal),
    .io_y_paa(entries_barrier_4_io_y_paa),
    .io_y_eff(entries_barrier_4_io_y_eff),
    .io_y_c(entries_barrier_4_io_y_c)
  );
  OptimizationBarrier entries_barrier_5 ( // @[package.scala 236:25]
    .io_x_ppn(entries_barrier_5_io_x_ppn),
    .io_x_u(entries_barrier_5_io_x_u),
    .io_x_ae(entries_barrier_5_io_x_ae),
    .io_x_sw(entries_barrier_5_io_x_sw),
    .io_x_sx(entries_barrier_5_io_x_sx),
    .io_x_sr(entries_barrier_5_io_x_sr),
    .io_x_pw(entries_barrier_5_io_x_pw),
    .io_x_px(entries_barrier_5_io_x_px),
    .io_x_pr(entries_barrier_5_io_x_pr),
    .io_x_ppp(entries_barrier_5_io_x_ppp),
    .io_x_pal(entries_barrier_5_io_x_pal),
    .io_x_paa(entries_barrier_5_io_x_paa),
    .io_x_eff(entries_barrier_5_io_x_eff),
    .io_x_c(entries_barrier_5_io_x_c),
    .io_y_ppn(entries_barrier_5_io_y_ppn),
    .io_y_u(entries_barrier_5_io_y_u),
    .io_y_ae(entries_barrier_5_io_y_ae),
    .io_y_sw(entries_barrier_5_io_y_sw),
    .io_y_sx(entries_barrier_5_io_y_sx),
    .io_y_sr(entries_barrier_5_io_y_sr),
    .io_y_pw(entries_barrier_5_io_y_pw),
    .io_y_px(entries_barrier_5_io_y_px),
    .io_y_pr(entries_barrier_5_io_y_pr),
    .io_y_ppp(entries_barrier_5_io_y_ppp),
    .io_y_pal(entries_barrier_5_io_y_pal),
    .io_y_paa(entries_barrier_5_io_y_paa),
    .io_y_eff(entries_barrier_5_io_y_eff),
    .io_y_c(entries_barrier_5_io_y_c)
  );
  OptimizationBarrier entries_barrier_6 ( // @[package.scala 236:25]
    .io_x_ppn(entries_barrier_6_io_x_ppn),
    .io_x_u(entries_barrier_6_io_x_u),
    .io_x_ae(entries_barrier_6_io_x_ae),
    .io_x_sw(entries_barrier_6_io_x_sw),
    .io_x_sx(entries_barrier_6_io_x_sx),
    .io_x_sr(entries_barrier_6_io_x_sr),
    .io_x_pw(entries_barrier_6_io_x_pw),
    .io_x_px(entries_barrier_6_io_x_px),
    .io_x_pr(entries_barrier_6_io_x_pr),
    .io_x_ppp(entries_barrier_6_io_x_ppp),
    .io_x_pal(entries_barrier_6_io_x_pal),
    .io_x_paa(entries_barrier_6_io_x_paa),
    .io_x_eff(entries_barrier_6_io_x_eff),
    .io_x_c(entries_barrier_6_io_x_c),
    .io_y_ppn(entries_barrier_6_io_y_ppn),
    .io_y_u(entries_barrier_6_io_y_u),
    .io_y_ae(entries_barrier_6_io_y_ae),
    .io_y_sw(entries_barrier_6_io_y_sw),
    .io_y_sx(entries_barrier_6_io_y_sx),
    .io_y_sr(entries_barrier_6_io_y_sr),
    .io_y_pw(entries_barrier_6_io_y_pw),
    .io_y_px(entries_barrier_6_io_y_px),
    .io_y_pr(entries_barrier_6_io_y_pr),
    .io_y_ppp(entries_barrier_6_io_y_ppp),
    .io_y_pal(entries_barrier_6_io_y_pal),
    .io_y_paa(entries_barrier_6_io_y_paa),
    .io_y_eff(entries_barrier_6_io_y_eff),
    .io_y_c(entries_barrier_6_io_y_c)
  );
  OptimizationBarrier entries_barrier_7 ( // @[package.scala 236:25]
    .io_x_ppn(entries_barrier_7_io_x_ppn),
    .io_x_u(entries_barrier_7_io_x_u),
    .io_x_ae(entries_barrier_7_io_x_ae),
    .io_x_sw(entries_barrier_7_io_x_sw),
    .io_x_sx(entries_barrier_7_io_x_sx),
    .io_x_sr(entries_barrier_7_io_x_sr),
    .io_x_pw(entries_barrier_7_io_x_pw),
    .io_x_px(entries_barrier_7_io_x_px),
    .io_x_pr(entries_barrier_7_io_x_pr),
    .io_x_ppp(entries_barrier_7_io_x_ppp),
    .io_x_pal(entries_barrier_7_io_x_pal),
    .io_x_paa(entries_barrier_7_io_x_paa),
    .io_x_eff(entries_barrier_7_io_x_eff),
    .io_x_c(entries_barrier_7_io_x_c),
    .io_y_ppn(entries_barrier_7_io_y_ppn),
    .io_y_u(entries_barrier_7_io_y_u),
    .io_y_ae(entries_barrier_7_io_y_ae),
    .io_y_sw(entries_barrier_7_io_y_sw),
    .io_y_sx(entries_barrier_7_io_y_sx),
    .io_y_sr(entries_barrier_7_io_y_sr),
    .io_y_pw(entries_barrier_7_io_y_pw),
    .io_y_px(entries_barrier_7_io_y_px),
    .io_y_pr(entries_barrier_7_io_y_pr),
    .io_y_ppp(entries_barrier_7_io_y_ppp),
    .io_y_pal(entries_barrier_7_io_y_pal),
    .io_y_paa(entries_barrier_7_io_y_paa),
    .io_y_eff(entries_barrier_7_io_y_eff),
    .io_y_c(entries_barrier_7_io_y_c)
  );
  OptimizationBarrier entries_barrier_8 ( // @[package.scala 236:25]
    .io_x_ppn(entries_barrier_8_io_x_ppn),
    .io_x_u(entries_barrier_8_io_x_u),
    .io_x_ae(entries_barrier_8_io_x_ae),
    .io_x_sw(entries_barrier_8_io_x_sw),
    .io_x_sx(entries_barrier_8_io_x_sx),
    .io_x_sr(entries_barrier_8_io_x_sr),
    .io_x_pw(entries_barrier_8_io_x_pw),
    .io_x_px(entries_barrier_8_io_x_px),
    .io_x_pr(entries_barrier_8_io_x_pr),
    .io_x_ppp(entries_barrier_8_io_x_ppp),
    .io_x_pal(entries_barrier_8_io_x_pal),
    .io_x_paa(entries_barrier_8_io_x_paa),
    .io_x_eff(entries_barrier_8_io_x_eff),
    .io_x_c(entries_barrier_8_io_x_c),
    .io_y_ppn(entries_barrier_8_io_y_ppn),
    .io_y_u(entries_barrier_8_io_y_u),
    .io_y_ae(entries_barrier_8_io_y_ae),
    .io_y_sw(entries_barrier_8_io_y_sw),
    .io_y_sx(entries_barrier_8_io_y_sx),
    .io_y_sr(entries_barrier_8_io_y_sr),
    .io_y_pw(entries_barrier_8_io_y_pw),
    .io_y_px(entries_barrier_8_io_y_px),
    .io_y_pr(entries_barrier_8_io_y_pr),
    .io_y_ppp(entries_barrier_8_io_y_ppp),
    .io_y_pal(entries_barrier_8_io_y_pal),
    .io_y_paa(entries_barrier_8_io_y_paa),
    .io_y_eff(entries_barrier_8_io_y_eff),
    .io_y_c(entries_barrier_8_io_y_c)
  );
  OptimizationBarrier entries_barrier_9 ( // @[package.scala 236:25]
    .io_x_ppn(entries_barrier_9_io_x_ppn),
    .io_x_u(entries_barrier_9_io_x_u),
    .io_x_ae(entries_barrier_9_io_x_ae),
    .io_x_sw(entries_barrier_9_io_x_sw),
    .io_x_sx(entries_barrier_9_io_x_sx),
    .io_x_sr(entries_barrier_9_io_x_sr),
    .io_x_pw(entries_barrier_9_io_x_pw),
    .io_x_px(entries_barrier_9_io_x_px),
    .io_x_pr(entries_barrier_9_io_x_pr),
    .io_x_ppp(entries_barrier_9_io_x_ppp),
    .io_x_pal(entries_barrier_9_io_x_pal),
    .io_x_paa(entries_barrier_9_io_x_paa),
    .io_x_eff(entries_barrier_9_io_x_eff),
    .io_x_c(entries_barrier_9_io_x_c),
    .io_y_ppn(entries_barrier_9_io_y_ppn),
    .io_y_u(entries_barrier_9_io_y_u),
    .io_y_ae(entries_barrier_9_io_y_ae),
    .io_y_sw(entries_barrier_9_io_y_sw),
    .io_y_sx(entries_barrier_9_io_y_sx),
    .io_y_sr(entries_barrier_9_io_y_sr),
    .io_y_pw(entries_barrier_9_io_y_pw),
    .io_y_px(entries_barrier_9_io_y_px),
    .io_y_pr(entries_barrier_9_io_y_pr),
    .io_y_ppp(entries_barrier_9_io_y_ppp),
    .io_y_pal(entries_barrier_9_io_y_pal),
    .io_y_paa(entries_barrier_9_io_y_paa),
    .io_y_eff(entries_barrier_9_io_y_eff),
    .io_y_c(entries_barrier_9_io_y_c)
  );
  OptimizationBarrier entries_barrier_10 ( // @[package.scala 236:25]
    .io_x_ppn(entries_barrier_10_io_x_ppn),
    .io_x_u(entries_barrier_10_io_x_u),
    .io_x_ae(entries_barrier_10_io_x_ae),
    .io_x_sw(entries_barrier_10_io_x_sw),
    .io_x_sx(entries_barrier_10_io_x_sx),
    .io_x_sr(entries_barrier_10_io_x_sr),
    .io_x_pw(entries_barrier_10_io_x_pw),
    .io_x_px(entries_barrier_10_io_x_px),
    .io_x_pr(entries_barrier_10_io_x_pr),
    .io_x_ppp(entries_barrier_10_io_x_ppp),
    .io_x_pal(entries_barrier_10_io_x_pal),
    .io_x_paa(entries_barrier_10_io_x_paa),
    .io_x_eff(entries_barrier_10_io_x_eff),
    .io_x_c(entries_barrier_10_io_x_c),
    .io_y_ppn(entries_barrier_10_io_y_ppn),
    .io_y_u(entries_barrier_10_io_y_u),
    .io_y_ae(entries_barrier_10_io_y_ae),
    .io_y_sw(entries_barrier_10_io_y_sw),
    .io_y_sx(entries_barrier_10_io_y_sx),
    .io_y_sr(entries_barrier_10_io_y_sr),
    .io_y_pw(entries_barrier_10_io_y_pw),
    .io_y_px(entries_barrier_10_io_y_px),
    .io_y_pr(entries_barrier_10_io_y_pr),
    .io_y_ppp(entries_barrier_10_io_y_ppp),
    .io_y_pal(entries_barrier_10_io_y_pal),
    .io_y_paa(entries_barrier_10_io_y_paa),
    .io_y_eff(entries_barrier_10_io_y_eff),
    .io_y_c(entries_barrier_10_io_y_c)
  );
  OptimizationBarrier entries_barrier_11 ( // @[package.scala 236:25]
    .io_x_ppn(entries_barrier_11_io_x_ppn),
    .io_x_u(entries_barrier_11_io_x_u),
    .io_x_ae(entries_barrier_11_io_x_ae),
    .io_x_sw(entries_barrier_11_io_x_sw),
    .io_x_sx(entries_barrier_11_io_x_sx),
    .io_x_sr(entries_barrier_11_io_x_sr),
    .io_x_pw(entries_barrier_11_io_x_pw),
    .io_x_px(entries_barrier_11_io_x_px),
    .io_x_pr(entries_barrier_11_io_x_pr),
    .io_x_ppp(entries_barrier_11_io_x_ppp),
    .io_x_pal(entries_barrier_11_io_x_pal),
    .io_x_paa(entries_barrier_11_io_x_paa),
    .io_x_eff(entries_barrier_11_io_x_eff),
    .io_x_c(entries_barrier_11_io_x_c),
    .io_y_ppn(entries_barrier_11_io_y_ppn),
    .io_y_u(entries_barrier_11_io_y_u),
    .io_y_ae(entries_barrier_11_io_y_ae),
    .io_y_sw(entries_barrier_11_io_y_sw),
    .io_y_sx(entries_barrier_11_io_y_sx),
    .io_y_sr(entries_barrier_11_io_y_sr),
    .io_y_pw(entries_barrier_11_io_y_pw),
    .io_y_px(entries_barrier_11_io_y_px),
    .io_y_pr(entries_barrier_11_io_y_pr),
    .io_y_ppp(entries_barrier_11_io_y_ppp),
    .io_y_pal(entries_barrier_11_io_y_pal),
    .io_y_paa(entries_barrier_11_io_y_paa),
    .io_y_eff(entries_barrier_11_io_y_eff),
    .io_y_c(entries_barrier_11_io_y_c)
  );
  OptimizationBarrier entries_barrier_12 ( // @[package.scala 236:25]
    .io_x_ppn(entries_barrier_12_io_x_ppn),
    .io_x_u(entries_barrier_12_io_x_u),
    .io_x_ae(entries_barrier_12_io_x_ae),
    .io_x_sw(entries_barrier_12_io_x_sw),
    .io_x_sx(entries_barrier_12_io_x_sx),
    .io_x_sr(entries_barrier_12_io_x_sr),
    .io_x_pw(entries_barrier_12_io_x_pw),
    .io_x_px(entries_barrier_12_io_x_px),
    .io_x_pr(entries_barrier_12_io_x_pr),
    .io_x_ppp(entries_barrier_12_io_x_ppp),
    .io_x_pal(entries_barrier_12_io_x_pal),
    .io_x_paa(entries_barrier_12_io_x_paa),
    .io_x_eff(entries_barrier_12_io_x_eff),
    .io_x_c(entries_barrier_12_io_x_c),
    .io_y_ppn(entries_barrier_12_io_y_ppn),
    .io_y_u(entries_barrier_12_io_y_u),
    .io_y_ae(entries_barrier_12_io_y_ae),
    .io_y_sw(entries_barrier_12_io_y_sw),
    .io_y_sx(entries_barrier_12_io_y_sx),
    .io_y_sr(entries_barrier_12_io_y_sr),
    .io_y_pw(entries_barrier_12_io_y_pw),
    .io_y_px(entries_barrier_12_io_y_px),
    .io_y_pr(entries_barrier_12_io_y_pr),
    .io_y_ppp(entries_barrier_12_io_y_ppp),
    .io_y_pal(entries_barrier_12_io_y_pal),
    .io_y_paa(entries_barrier_12_io_y_paa),
    .io_y_eff(entries_barrier_12_io_y_eff),
    .io_y_c(entries_barrier_12_io_y_c)
  );
  OptimizationBarrier normal_entries_barrier ( // @[package.scala 236:25]
    .io_x_ppn(normal_entries_barrier_io_x_ppn),
    .io_x_u(normal_entries_barrier_io_x_u),
    .io_x_ae(normal_entries_barrier_io_x_ae),
    .io_x_sw(normal_entries_barrier_io_x_sw),
    .io_x_sx(normal_entries_barrier_io_x_sx),
    .io_x_sr(normal_entries_barrier_io_x_sr),
    .io_x_pw(normal_entries_barrier_io_x_pw),
    .io_x_px(normal_entries_barrier_io_x_px),
    .io_x_pr(normal_entries_barrier_io_x_pr),
    .io_x_ppp(normal_entries_barrier_io_x_ppp),
    .io_x_pal(normal_entries_barrier_io_x_pal),
    .io_x_paa(normal_entries_barrier_io_x_paa),
    .io_x_eff(normal_entries_barrier_io_x_eff),
    .io_x_c(normal_entries_barrier_io_x_c),
    .io_y_ppn(normal_entries_barrier_io_y_ppn),
    .io_y_u(normal_entries_barrier_io_y_u),
    .io_y_ae(normal_entries_barrier_io_y_ae),
    .io_y_sw(normal_entries_barrier_io_y_sw),
    .io_y_sx(normal_entries_barrier_io_y_sx),
    .io_y_sr(normal_entries_barrier_io_y_sr),
    .io_y_pw(normal_entries_barrier_io_y_pw),
    .io_y_px(normal_entries_barrier_io_y_px),
    .io_y_pr(normal_entries_barrier_io_y_pr),
    .io_y_ppp(normal_entries_barrier_io_y_ppp),
    .io_y_pal(normal_entries_barrier_io_y_pal),
    .io_y_paa(normal_entries_barrier_io_y_paa),
    .io_y_eff(normal_entries_barrier_io_y_eff),
    .io_y_c(normal_entries_barrier_io_y_c)
  );
  OptimizationBarrier normal_entries_barrier_1 ( // @[package.scala 236:25]
    .io_x_ppn(normal_entries_barrier_1_io_x_ppn),
    .io_x_u(normal_entries_barrier_1_io_x_u),
    .io_x_ae(normal_entries_barrier_1_io_x_ae),
    .io_x_sw(normal_entries_barrier_1_io_x_sw),
    .io_x_sx(normal_entries_barrier_1_io_x_sx),
    .io_x_sr(normal_entries_barrier_1_io_x_sr),
    .io_x_pw(normal_entries_barrier_1_io_x_pw),
    .io_x_px(normal_entries_barrier_1_io_x_px),
    .io_x_pr(normal_entries_barrier_1_io_x_pr),
    .io_x_ppp(normal_entries_barrier_1_io_x_ppp),
    .io_x_pal(normal_entries_barrier_1_io_x_pal),
    .io_x_paa(normal_entries_barrier_1_io_x_paa),
    .io_x_eff(normal_entries_barrier_1_io_x_eff),
    .io_x_c(normal_entries_barrier_1_io_x_c),
    .io_y_ppn(normal_entries_barrier_1_io_y_ppn),
    .io_y_u(normal_entries_barrier_1_io_y_u),
    .io_y_ae(normal_entries_barrier_1_io_y_ae),
    .io_y_sw(normal_entries_barrier_1_io_y_sw),
    .io_y_sx(normal_entries_barrier_1_io_y_sx),
    .io_y_sr(normal_entries_barrier_1_io_y_sr),
    .io_y_pw(normal_entries_barrier_1_io_y_pw),
    .io_y_px(normal_entries_barrier_1_io_y_px),
    .io_y_pr(normal_entries_barrier_1_io_y_pr),
    .io_y_ppp(normal_entries_barrier_1_io_y_ppp),
    .io_y_pal(normal_entries_barrier_1_io_y_pal),
    .io_y_paa(normal_entries_barrier_1_io_y_paa),
    .io_y_eff(normal_entries_barrier_1_io_y_eff),
    .io_y_c(normal_entries_barrier_1_io_y_c)
  );
  OptimizationBarrier normal_entries_barrier_2 ( // @[package.scala 236:25]
    .io_x_ppn(normal_entries_barrier_2_io_x_ppn),
    .io_x_u(normal_entries_barrier_2_io_x_u),
    .io_x_ae(normal_entries_barrier_2_io_x_ae),
    .io_x_sw(normal_entries_barrier_2_io_x_sw),
    .io_x_sx(normal_entries_barrier_2_io_x_sx),
    .io_x_sr(normal_entries_barrier_2_io_x_sr),
    .io_x_pw(normal_entries_barrier_2_io_x_pw),
    .io_x_px(normal_entries_barrier_2_io_x_px),
    .io_x_pr(normal_entries_barrier_2_io_x_pr),
    .io_x_ppp(normal_entries_barrier_2_io_x_ppp),
    .io_x_pal(normal_entries_barrier_2_io_x_pal),
    .io_x_paa(normal_entries_barrier_2_io_x_paa),
    .io_x_eff(normal_entries_barrier_2_io_x_eff),
    .io_x_c(normal_entries_barrier_2_io_x_c),
    .io_y_ppn(normal_entries_barrier_2_io_y_ppn),
    .io_y_u(normal_entries_barrier_2_io_y_u),
    .io_y_ae(normal_entries_barrier_2_io_y_ae),
    .io_y_sw(normal_entries_barrier_2_io_y_sw),
    .io_y_sx(normal_entries_barrier_2_io_y_sx),
    .io_y_sr(normal_entries_barrier_2_io_y_sr),
    .io_y_pw(normal_entries_barrier_2_io_y_pw),
    .io_y_px(normal_entries_barrier_2_io_y_px),
    .io_y_pr(normal_entries_barrier_2_io_y_pr),
    .io_y_ppp(normal_entries_barrier_2_io_y_ppp),
    .io_y_pal(normal_entries_barrier_2_io_y_pal),
    .io_y_paa(normal_entries_barrier_2_io_y_paa),
    .io_y_eff(normal_entries_barrier_2_io_y_eff),
    .io_y_c(normal_entries_barrier_2_io_y_c)
  );
  OptimizationBarrier normal_entries_barrier_3 ( // @[package.scala 236:25]
    .io_x_ppn(normal_entries_barrier_3_io_x_ppn),
    .io_x_u(normal_entries_barrier_3_io_x_u),
    .io_x_ae(normal_entries_barrier_3_io_x_ae),
    .io_x_sw(normal_entries_barrier_3_io_x_sw),
    .io_x_sx(normal_entries_barrier_3_io_x_sx),
    .io_x_sr(normal_entries_barrier_3_io_x_sr),
    .io_x_pw(normal_entries_barrier_3_io_x_pw),
    .io_x_px(normal_entries_barrier_3_io_x_px),
    .io_x_pr(normal_entries_barrier_3_io_x_pr),
    .io_x_ppp(normal_entries_barrier_3_io_x_ppp),
    .io_x_pal(normal_entries_barrier_3_io_x_pal),
    .io_x_paa(normal_entries_barrier_3_io_x_paa),
    .io_x_eff(normal_entries_barrier_3_io_x_eff),
    .io_x_c(normal_entries_barrier_3_io_x_c),
    .io_y_ppn(normal_entries_barrier_3_io_y_ppn),
    .io_y_u(normal_entries_barrier_3_io_y_u),
    .io_y_ae(normal_entries_barrier_3_io_y_ae),
    .io_y_sw(normal_entries_barrier_3_io_y_sw),
    .io_y_sx(normal_entries_barrier_3_io_y_sx),
    .io_y_sr(normal_entries_barrier_3_io_y_sr),
    .io_y_pw(normal_entries_barrier_3_io_y_pw),
    .io_y_px(normal_entries_barrier_3_io_y_px),
    .io_y_pr(normal_entries_barrier_3_io_y_pr),
    .io_y_ppp(normal_entries_barrier_3_io_y_ppp),
    .io_y_pal(normal_entries_barrier_3_io_y_pal),
    .io_y_paa(normal_entries_barrier_3_io_y_paa),
    .io_y_eff(normal_entries_barrier_3_io_y_eff),
    .io_y_c(normal_entries_barrier_3_io_y_c)
  );
  OptimizationBarrier normal_entries_barrier_4 ( // @[package.scala 236:25]
    .io_x_ppn(normal_entries_barrier_4_io_x_ppn),
    .io_x_u(normal_entries_barrier_4_io_x_u),
    .io_x_ae(normal_entries_barrier_4_io_x_ae),
    .io_x_sw(normal_entries_barrier_4_io_x_sw),
    .io_x_sx(normal_entries_barrier_4_io_x_sx),
    .io_x_sr(normal_entries_barrier_4_io_x_sr),
    .io_x_pw(normal_entries_barrier_4_io_x_pw),
    .io_x_px(normal_entries_barrier_4_io_x_px),
    .io_x_pr(normal_entries_barrier_4_io_x_pr),
    .io_x_ppp(normal_entries_barrier_4_io_x_ppp),
    .io_x_pal(normal_entries_barrier_4_io_x_pal),
    .io_x_paa(normal_entries_barrier_4_io_x_paa),
    .io_x_eff(normal_entries_barrier_4_io_x_eff),
    .io_x_c(normal_entries_barrier_4_io_x_c),
    .io_y_ppn(normal_entries_barrier_4_io_y_ppn),
    .io_y_u(normal_entries_barrier_4_io_y_u),
    .io_y_ae(normal_entries_barrier_4_io_y_ae),
    .io_y_sw(normal_entries_barrier_4_io_y_sw),
    .io_y_sx(normal_entries_barrier_4_io_y_sx),
    .io_y_sr(normal_entries_barrier_4_io_y_sr),
    .io_y_pw(normal_entries_barrier_4_io_y_pw),
    .io_y_px(normal_entries_barrier_4_io_y_px),
    .io_y_pr(normal_entries_barrier_4_io_y_pr),
    .io_y_ppp(normal_entries_barrier_4_io_y_ppp),
    .io_y_pal(normal_entries_barrier_4_io_y_pal),
    .io_y_paa(normal_entries_barrier_4_io_y_paa),
    .io_y_eff(normal_entries_barrier_4_io_y_eff),
    .io_y_c(normal_entries_barrier_4_io_y_c)
  );
  OptimizationBarrier normal_entries_barrier_5 ( // @[package.scala 236:25]
    .io_x_ppn(normal_entries_barrier_5_io_x_ppn),
    .io_x_u(normal_entries_barrier_5_io_x_u),
    .io_x_ae(normal_entries_barrier_5_io_x_ae),
    .io_x_sw(normal_entries_barrier_5_io_x_sw),
    .io_x_sx(normal_entries_barrier_5_io_x_sx),
    .io_x_sr(normal_entries_barrier_5_io_x_sr),
    .io_x_pw(normal_entries_barrier_5_io_x_pw),
    .io_x_px(normal_entries_barrier_5_io_x_px),
    .io_x_pr(normal_entries_barrier_5_io_x_pr),
    .io_x_ppp(normal_entries_barrier_5_io_x_ppp),
    .io_x_pal(normal_entries_barrier_5_io_x_pal),
    .io_x_paa(normal_entries_barrier_5_io_x_paa),
    .io_x_eff(normal_entries_barrier_5_io_x_eff),
    .io_x_c(normal_entries_barrier_5_io_x_c),
    .io_y_ppn(normal_entries_barrier_5_io_y_ppn),
    .io_y_u(normal_entries_barrier_5_io_y_u),
    .io_y_ae(normal_entries_barrier_5_io_y_ae),
    .io_y_sw(normal_entries_barrier_5_io_y_sw),
    .io_y_sx(normal_entries_barrier_5_io_y_sx),
    .io_y_sr(normal_entries_barrier_5_io_y_sr),
    .io_y_pw(normal_entries_barrier_5_io_y_pw),
    .io_y_px(normal_entries_barrier_5_io_y_px),
    .io_y_pr(normal_entries_barrier_5_io_y_pr),
    .io_y_ppp(normal_entries_barrier_5_io_y_ppp),
    .io_y_pal(normal_entries_barrier_5_io_y_pal),
    .io_y_paa(normal_entries_barrier_5_io_y_paa),
    .io_y_eff(normal_entries_barrier_5_io_y_eff),
    .io_y_c(normal_entries_barrier_5_io_y_c)
  );
  OptimizationBarrier normal_entries_barrier_6 ( // @[package.scala 236:25]
    .io_x_ppn(normal_entries_barrier_6_io_x_ppn),
    .io_x_u(normal_entries_barrier_6_io_x_u),
    .io_x_ae(normal_entries_barrier_6_io_x_ae),
    .io_x_sw(normal_entries_barrier_6_io_x_sw),
    .io_x_sx(normal_entries_barrier_6_io_x_sx),
    .io_x_sr(normal_entries_barrier_6_io_x_sr),
    .io_x_pw(normal_entries_barrier_6_io_x_pw),
    .io_x_px(normal_entries_barrier_6_io_x_px),
    .io_x_pr(normal_entries_barrier_6_io_x_pr),
    .io_x_ppp(normal_entries_barrier_6_io_x_ppp),
    .io_x_pal(normal_entries_barrier_6_io_x_pal),
    .io_x_paa(normal_entries_barrier_6_io_x_paa),
    .io_x_eff(normal_entries_barrier_6_io_x_eff),
    .io_x_c(normal_entries_barrier_6_io_x_c),
    .io_y_ppn(normal_entries_barrier_6_io_y_ppn),
    .io_y_u(normal_entries_barrier_6_io_y_u),
    .io_y_ae(normal_entries_barrier_6_io_y_ae),
    .io_y_sw(normal_entries_barrier_6_io_y_sw),
    .io_y_sx(normal_entries_barrier_6_io_y_sx),
    .io_y_sr(normal_entries_barrier_6_io_y_sr),
    .io_y_pw(normal_entries_barrier_6_io_y_pw),
    .io_y_px(normal_entries_barrier_6_io_y_px),
    .io_y_pr(normal_entries_barrier_6_io_y_pr),
    .io_y_ppp(normal_entries_barrier_6_io_y_ppp),
    .io_y_pal(normal_entries_barrier_6_io_y_pal),
    .io_y_paa(normal_entries_barrier_6_io_y_paa),
    .io_y_eff(normal_entries_barrier_6_io_y_eff),
    .io_y_c(normal_entries_barrier_6_io_y_c)
  );
  OptimizationBarrier normal_entries_barrier_7 ( // @[package.scala 236:25]
    .io_x_ppn(normal_entries_barrier_7_io_x_ppn),
    .io_x_u(normal_entries_barrier_7_io_x_u),
    .io_x_ae(normal_entries_barrier_7_io_x_ae),
    .io_x_sw(normal_entries_barrier_7_io_x_sw),
    .io_x_sx(normal_entries_barrier_7_io_x_sx),
    .io_x_sr(normal_entries_barrier_7_io_x_sr),
    .io_x_pw(normal_entries_barrier_7_io_x_pw),
    .io_x_px(normal_entries_barrier_7_io_x_px),
    .io_x_pr(normal_entries_barrier_7_io_x_pr),
    .io_x_ppp(normal_entries_barrier_7_io_x_ppp),
    .io_x_pal(normal_entries_barrier_7_io_x_pal),
    .io_x_paa(normal_entries_barrier_7_io_x_paa),
    .io_x_eff(normal_entries_barrier_7_io_x_eff),
    .io_x_c(normal_entries_barrier_7_io_x_c),
    .io_y_ppn(normal_entries_barrier_7_io_y_ppn),
    .io_y_u(normal_entries_barrier_7_io_y_u),
    .io_y_ae(normal_entries_barrier_7_io_y_ae),
    .io_y_sw(normal_entries_barrier_7_io_y_sw),
    .io_y_sx(normal_entries_barrier_7_io_y_sx),
    .io_y_sr(normal_entries_barrier_7_io_y_sr),
    .io_y_pw(normal_entries_barrier_7_io_y_pw),
    .io_y_px(normal_entries_barrier_7_io_y_px),
    .io_y_pr(normal_entries_barrier_7_io_y_pr),
    .io_y_ppp(normal_entries_barrier_7_io_y_ppp),
    .io_y_pal(normal_entries_barrier_7_io_y_pal),
    .io_y_paa(normal_entries_barrier_7_io_y_paa),
    .io_y_eff(normal_entries_barrier_7_io_y_eff),
    .io_y_c(normal_entries_barrier_7_io_y_c)
  );
  OptimizationBarrier normal_entries_barrier_8 ( // @[package.scala 236:25]
    .io_x_ppn(normal_entries_barrier_8_io_x_ppn),
    .io_x_u(normal_entries_barrier_8_io_x_u),
    .io_x_ae(normal_entries_barrier_8_io_x_ae),
    .io_x_sw(normal_entries_barrier_8_io_x_sw),
    .io_x_sx(normal_entries_barrier_8_io_x_sx),
    .io_x_sr(normal_entries_barrier_8_io_x_sr),
    .io_x_pw(normal_entries_barrier_8_io_x_pw),
    .io_x_px(normal_entries_barrier_8_io_x_px),
    .io_x_pr(normal_entries_barrier_8_io_x_pr),
    .io_x_ppp(normal_entries_barrier_8_io_x_ppp),
    .io_x_pal(normal_entries_barrier_8_io_x_pal),
    .io_x_paa(normal_entries_barrier_8_io_x_paa),
    .io_x_eff(normal_entries_barrier_8_io_x_eff),
    .io_x_c(normal_entries_barrier_8_io_x_c),
    .io_y_ppn(normal_entries_barrier_8_io_y_ppn),
    .io_y_u(normal_entries_barrier_8_io_y_u),
    .io_y_ae(normal_entries_barrier_8_io_y_ae),
    .io_y_sw(normal_entries_barrier_8_io_y_sw),
    .io_y_sx(normal_entries_barrier_8_io_y_sx),
    .io_y_sr(normal_entries_barrier_8_io_y_sr),
    .io_y_pw(normal_entries_barrier_8_io_y_pw),
    .io_y_px(normal_entries_barrier_8_io_y_px),
    .io_y_pr(normal_entries_barrier_8_io_y_pr),
    .io_y_ppp(normal_entries_barrier_8_io_y_ppp),
    .io_y_pal(normal_entries_barrier_8_io_y_pal),
    .io_y_paa(normal_entries_barrier_8_io_y_paa),
    .io_y_eff(normal_entries_barrier_8_io_y_eff),
    .io_y_c(normal_entries_barrier_8_io_y_c)
  );
  OptimizationBarrier normal_entries_barrier_9 ( // @[package.scala 236:25]
    .io_x_ppn(normal_entries_barrier_9_io_x_ppn),
    .io_x_u(normal_entries_barrier_9_io_x_u),
    .io_x_ae(normal_entries_barrier_9_io_x_ae),
    .io_x_sw(normal_entries_barrier_9_io_x_sw),
    .io_x_sx(normal_entries_barrier_9_io_x_sx),
    .io_x_sr(normal_entries_barrier_9_io_x_sr),
    .io_x_pw(normal_entries_barrier_9_io_x_pw),
    .io_x_px(normal_entries_barrier_9_io_x_px),
    .io_x_pr(normal_entries_barrier_9_io_x_pr),
    .io_x_ppp(normal_entries_barrier_9_io_x_ppp),
    .io_x_pal(normal_entries_barrier_9_io_x_pal),
    .io_x_paa(normal_entries_barrier_9_io_x_paa),
    .io_x_eff(normal_entries_barrier_9_io_x_eff),
    .io_x_c(normal_entries_barrier_9_io_x_c),
    .io_y_ppn(normal_entries_barrier_9_io_y_ppn),
    .io_y_u(normal_entries_barrier_9_io_y_u),
    .io_y_ae(normal_entries_barrier_9_io_y_ae),
    .io_y_sw(normal_entries_barrier_9_io_y_sw),
    .io_y_sx(normal_entries_barrier_9_io_y_sx),
    .io_y_sr(normal_entries_barrier_9_io_y_sr),
    .io_y_pw(normal_entries_barrier_9_io_y_pw),
    .io_y_px(normal_entries_barrier_9_io_y_px),
    .io_y_pr(normal_entries_barrier_9_io_y_pr),
    .io_y_ppp(normal_entries_barrier_9_io_y_ppp),
    .io_y_pal(normal_entries_barrier_9_io_y_pal),
    .io_y_paa(normal_entries_barrier_9_io_y_paa),
    .io_y_eff(normal_entries_barrier_9_io_y_eff),
    .io_y_c(normal_entries_barrier_9_io_y_c)
  );
  OptimizationBarrier normal_entries_barrier_10 ( // @[package.scala 236:25]
    .io_x_ppn(normal_entries_barrier_10_io_x_ppn),
    .io_x_u(normal_entries_barrier_10_io_x_u),
    .io_x_ae(normal_entries_barrier_10_io_x_ae),
    .io_x_sw(normal_entries_barrier_10_io_x_sw),
    .io_x_sx(normal_entries_barrier_10_io_x_sx),
    .io_x_sr(normal_entries_barrier_10_io_x_sr),
    .io_x_pw(normal_entries_barrier_10_io_x_pw),
    .io_x_px(normal_entries_barrier_10_io_x_px),
    .io_x_pr(normal_entries_barrier_10_io_x_pr),
    .io_x_ppp(normal_entries_barrier_10_io_x_ppp),
    .io_x_pal(normal_entries_barrier_10_io_x_pal),
    .io_x_paa(normal_entries_barrier_10_io_x_paa),
    .io_x_eff(normal_entries_barrier_10_io_x_eff),
    .io_x_c(normal_entries_barrier_10_io_x_c),
    .io_y_ppn(normal_entries_barrier_10_io_y_ppn),
    .io_y_u(normal_entries_barrier_10_io_y_u),
    .io_y_ae(normal_entries_barrier_10_io_y_ae),
    .io_y_sw(normal_entries_barrier_10_io_y_sw),
    .io_y_sx(normal_entries_barrier_10_io_y_sx),
    .io_y_sr(normal_entries_barrier_10_io_y_sr),
    .io_y_pw(normal_entries_barrier_10_io_y_pw),
    .io_y_px(normal_entries_barrier_10_io_y_px),
    .io_y_pr(normal_entries_barrier_10_io_y_pr),
    .io_y_ppp(normal_entries_barrier_10_io_y_ppp),
    .io_y_pal(normal_entries_barrier_10_io_y_pal),
    .io_y_paa(normal_entries_barrier_10_io_y_paa),
    .io_y_eff(normal_entries_barrier_10_io_y_eff),
    .io_y_c(normal_entries_barrier_10_io_y_c)
  );
  OptimizationBarrier normal_entries_barrier_11 ( // @[package.scala 236:25]
    .io_x_ppn(normal_entries_barrier_11_io_x_ppn),
    .io_x_u(normal_entries_barrier_11_io_x_u),
    .io_x_ae(normal_entries_barrier_11_io_x_ae),
    .io_x_sw(normal_entries_barrier_11_io_x_sw),
    .io_x_sx(normal_entries_barrier_11_io_x_sx),
    .io_x_sr(normal_entries_barrier_11_io_x_sr),
    .io_x_pw(normal_entries_barrier_11_io_x_pw),
    .io_x_px(normal_entries_barrier_11_io_x_px),
    .io_x_pr(normal_entries_barrier_11_io_x_pr),
    .io_x_ppp(normal_entries_barrier_11_io_x_ppp),
    .io_x_pal(normal_entries_barrier_11_io_x_pal),
    .io_x_paa(normal_entries_barrier_11_io_x_paa),
    .io_x_eff(normal_entries_barrier_11_io_x_eff),
    .io_x_c(normal_entries_barrier_11_io_x_c),
    .io_y_ppn(normal_entries_barrier_11_io_y_ppn),
    .io_y_u(normal_entries_barrier_11_io_y_u),
    .io_y_ae(normal_entries_barrier_11_io_y_ae),
    .io_y_sw(normal_entries_barrier_11_io_y_sw),
    .io_y_sx(normal_entries_barrier_11_io_y_sx),
    .io_y_sr(normal_entries_barrier_11_io_y_sr),
    .io_y_pw(normal_entries_barrier_11_io_y_pw),
    .io_y_px(normal_entries_barrier_11_io_y_px),
    .io_y_pr(normal_entries_barrier_11_io_y_pr),
    .io_y_ppp(normal_entries_barrier_11_io_y_ppp),
    .io_y_pal(normal_entries_barrier_11_io_y_pal),
    .io_y_paa(normal_entries_barrier_11_io_y_paa),
    .io_y_eff(normal_entries_barrier_11_io_y_eff),
    .io_y_c(normal_entries_barrier_11_io_y_c)
  );
  assign io_req_ready = state == 2'h0; // @[TLB.scala 337:25]
  assign io_resp_miss = (io_ptw_resp_valid | tlb_miss) | multipleHits; // @[TLB.scala 350:41]
  assign io_resp_paddr = {ppn,mpu_physaddr_left}; // @[Cat.scala 29:58]
  assign io_resp_pf_inst = bad_va | (|_io_resp_pf_inst_T); // @[TLB.scala 340:29]
  assign io_resp_ae_inst = |_io_resp_ae_inst_T_1; // @[TLB.scala 343:41]
  assign io_resp_cacheable = |_io_resp_cacheable_T; // @[TLB.scala 347:41]
  assign io_ptw_req_valid = state == 2'h1; // @[TLB.scala 353:29]
  assign io_ptw_req_bits_valid = ~io_kill; // @[TLB.scala 354:28]
  assign io_ptw_req_bits_bits_addr = r_refill_tag; // @[TLB.scala 355:29]
  assign mpu_ppn_data_barrier_io_x_ppn = special_entry_data_0[34:15]; // @[TLB.scala 86:77]
  assign mpu_ppn_data_barrier_io_x_u = special_entry_data_0[14]; // @[TLB.scala 86:77]
  assign mpu_ppn_data_barrier_io_x_ae = special_entry_data_0[12]; // @[TLB.scala 86:77]
  assign mpu_ppn_data_barrier_io_x_sw = special_entry_data_0[11]; // @[TLB.scala 86:77]
  assign mpu_ppn_data_barrier_io_x_sx = special_entry_data_0[10]; // @[TLB.scala 86:77]
  assign mpu_ppn_data_barrier_io_x_sr = special_entry_data_0[9]; // @[TLB.scala 86:77]
  assign mpu_ppn_data_barrier_io_x_pw = special_entry_data_0[8]; // @[TLB.scala 86:77]
  assign mpu_ppn_data_barrier_io_x_px = special_entry_data_0[7]; // @[TLB.scala 86:77]
  assign mpu_ppn_data_barrier_io_x_pr = special_entry_data_0[6]; // @[TLB.scala 86:77]
  assign mpu_ppn_data_barrier_io_x_ppp = special_entry_data_0[5]; // @[TLB.scala 86:77]
  assign mpu_ppn_data_barrier_io_x_pal = special_entry_data_0[4]; // @[TLB.scala 86:77]
  assign mpu_ppn_data_barrier_io_x_paa = special_entry_data_0[3]; // @[TLB.scala 86:77]
  assign mpu_ppn_data_barrier_io_x_eff = special_entry_data_0[2]; // @[TLB.scala 86:77]
  assign mpu_ppn_data_barrier_io_x_c = special_entry_data_0[1]; // @[TLB.scala 86:77]
  assign pmp_io_prv = mpu_priv[1:0]; // @[TLB.scala 194:14]
  assign pmp_io_pmp_0_cfg_l = io_ptw_pmp_0_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_0_cfg_a = io_ptw_pmp_0_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_0_cfg_x = io_ptw_pmp_0_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_0_cfg_w = io_ptw_pmp_0_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_0_cfg_r = io_ptw_pmp_0_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_0_addr = io_ptw_pmp_0_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_0_mask = io_ptw_pmp_0_mask; // @[TLB.scala 193:14]
  assign pmp_io_pmp_1_cfg_l = io_ptw_pmp_1_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_1_cfg_a = io_ptw_pmp_1_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_1_cfg_x = io_ptw_pmp_1_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_1_cfg_w = io_ptw_pmp_1_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_1_cfg_r = io_ptw_pmp_1_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_1_addr = io_ptw_pmp_1_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_1_mask = io_ptw_pmp_1_mask; // @[TLB.scala 193:14]
  assign pmp_io_pmp_2_cfg_l = io_ptw_pmp_2_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_2_cfg_a = io_ptw_pmp_2_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_2_cfg_x = io_ptw_pmp_2_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_2_cfg_w = io_ptw_pmp_2_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_2_cfg_r = io_ptw_pmp_2_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_2_addr = io_ptw_pmp_2_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_2_mask = io_ptw_pmp_2_mask; // @[TLB.scala 193:14]
  assign pmp_io_pmp_3_cfg_l = io_ptw_pmp_3_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_3_cfg_a = io_ptw_pmp_3_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_3_cfg_x = io_ptw_pmp_3_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_3_cfg_w = io_ptw_pmp_3_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_3_cfg_r = io_ptw_pmp_3_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_3_addr = io_ptw_pmp_3_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_3_mask = io_ptw_pmp_3_mask; // @[TLB.scala 193:14]
  assign pmp_io_pmp_4_cfg_l = io_ptw_pmp_4_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_4_cfg_a = io_ptw_pmp_4_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_4_cfg_x = io_ptw_pmp_4_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_4_cfg_w = io_ptw_pmp_4_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_4_cfg_r = io_ptw_pmp_4_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_4_addr = io_ptw_pmp_4_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_4_mask = io_ptw_pmp_4_mask; // @[TLB.scala 193:14]
  assign pmp_io_pmp_5_cfg_l = io_ptw_pmp_5_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_5_cfg_a = io_ptw_pmp_5_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_5_cfg_x = io_ptw_pmp_5_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_5_cfg_w = io_ptw_pmp_5_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_5_cfg_r = io_ptw_pmp_5_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_5_addr = io_ptw_pmp_5_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_5_mask = io_ptw_pmp_5_mask; // @[TLB.scala 193:14]
  assign pmp_io_pmp_6_cfg_l = io_ptw_pmp_6_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_6_cfg_a = io_ptw_pmp_6_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_6_cfg_x = io_ptw_pmp_6_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_6_cfg_w = io_ptw_pmp_6_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_6_cfg_r = io_ptw_pmp_6_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_6_addr = io_ptw_pmp_6_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_6_mask = io_ptw_pmp_6_mask; // @[TLB.scala 193:14]
  assign pmp_io_pmp_7_cfg_l = io_ptw_pmp_7_cfg_l; // @[TLB.scala 193:14]
  assign pmp_io_pmp_7_cfg_a = io_ptw_pmp_7_cfg_a; // @[TLB.scala 193:14]
  assign pmp_io_pmp_7_cfg_x = io_ptw_pmp_7_cfg_x; // @[TLB.scala 193:14]
  assign pmp_io_pmp_7_cfg_w = io_ptw_pmp_7_cfg_w; // @[TLB.scala 193:14]
  assign pmp_io_pmp_7_cfg_r = io_ptw_pmp_7_cfg_r; // @[TLB.scala 193:14]
  assign pmp_io_pmp_7_addr = io_ptw_pmp_7_addr; // @[TLB.scala 193:14]
  assign pmp_io_pmp_7_mask = io_ptw_pmp_7_mask; // @[TLB.scala 193:14]
  assign pmp_io_addr = mpu_physaddr[31:0]; // @[TLB.scala 191:15]
  assign ppn_data_barrier_io_x_ppn = _GEN_35[34:15]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_io_x_u = _GEN_35[14]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_io_x_ae = _GEN_35[12]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_io_x_sw = _GEN_35[11]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_io_x_sx = _GEN_35[10]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_io_x_sr = _GEN_35[9]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_io_x_pw = _GEN_35[8]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_io_x_px = _GEN_35[7]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_io_x_pr = _GEN_35[6]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_io_x_ppp = _GEN_35[5]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_io_x_pal = _GEN_35[4]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_io_x_paa = _GEN_35[3]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_io_x_eff = _GEN_35[2]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_io_x_c = _GEN_35[1]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_1_io_x_ppn = _GEN_39[34:15]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_1_io_x_u = _GEN_39[14]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_1_io_x_ae = _GEN_39[12]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_1_io_x_sw = _GEN_39[11]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_1_io_x_sx = _GEN_39[10]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_1_io_x_sr = _GEN_39[9]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_1_io_x_pw = _GEN_39[8]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_1_io_x_px = _GEN_39[7]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_1_io_x_pr = _GEN_39[6]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_1_io_x_ppp = _GEN_39[5]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_1_io_x_pal = _GEN_39[4]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_1_io_x_paa = _GEN_39[3]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_1_io_x_eff = _GEN_39[2]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_1_io_x_c = _GEN_39[1]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_2_io_x_ppn = _GEN_43[34:15]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_2_io_x_u = _GEN_43[14]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_2_io_x_ae = _GEN_43[12]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_2_io_x_sw = _GEN_43[11]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_2_io_x_sx = _GEN_43[10]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_2_io_x_sr = _GEN_43[9]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_2_io_x_pw = _GEN_43[8]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_2_io_x_px = _GEN_43[7]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_2_io_x_pr = _GEN_43[6]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_2_io_x_ppp = _GEN_43[5]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_2_io_x_pal = _GEN_43[4]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_2_io_x_paa = _GEN_43[3]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_2_io_x_eff = _GEN_43[2]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_2_io_x_c = _GEN_43[1]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_3_io_x_ppn = _GEN_47[34:15]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_3_io_x_u = _GEN_47[14]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_3_io_x_ae = _GEN_47[12]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_3_io_x_sw = _GEN_47[11]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_3_io_x_sx = _GEN_47[10]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_3_io_x_sr = _GEN_47[9]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_3_io_x_pw = _GEN_47[8]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_3_io_x_px = _GEN_47[7]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_3_io_x_pr = _GEN_47[6]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_3_io_x_ppp = _GEN_47[5]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_3_io_x_pal = _GEN_47[4]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_3_io_x_paa = _GEN_47[3]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_3_io_x_eff = _GEN_47[2]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_3_io_x_c = _GEN_47[1]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_4_io_x_ppn = _GEN_51[34:15]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_4_io_x_u = _GEN_51[14]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_4_io_x_ae = _GEN_51[12]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_4_io_x_sw = _GEN_51[11]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_4_io_x_sx = _GEN_51[10]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_4_io_x_sr = _GEN_51[9]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_4_io_x_pw = _GEN_51[8]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_4_io_x_px = _GEN_51[7]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_4_io_x_pr = _GEN_51[6]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_4_io_x_ppp = _GEN_51[5]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_4_io_x_pal = _GEN_51[4]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_4_io_x_paa = _GEN_51[3]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_4_io_x_eff = _GEN_51[2]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_4_io_x_c = _GEN_51[1]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_5_io_x_ppn = _GEN_55[34:15]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_5_io_x_u = _GEN_55[14]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_5_io_x_ae = _GEN_55[12]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_5_io_x_sw = _GEN_55[11]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_5_io_x_sx = _GEN_55[10]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_5_io_x_sr = _GEN_55[9]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_5_io_x_pw = _GEN_55[8]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_5_io_x_px = _GEN_55[7]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_5_io_x_pr = _GEN_55[6]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_5_io_x_ppp = _GEN_55[5]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_5_io_x_pal = _GEN_55[4]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_5_io_x_paa = _GEN_55[3]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_5_io_x_eff = _GEN_55[2]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_5_io_x_c = _GEN_55[1]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_6_io_x_ppn = _GEN_59[34:15]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_6_io_x_u = _GEN_59[14]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_6_io_x_ae = _GEN_59[12]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_6_io_x_sw = _GEN_59[11]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_6_io_x_sx = _GEN_59[10]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_6_io_x_sr = _GEN_59[9]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_6_io_x_pw = _GEN_59[8]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_6_io_x_px = _GEN_59[7]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_6_io_x_pr = _GEN_59[6]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_6_io_x_ppp = _GEN_59[5]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_6_io_x_pal = _GEN_59[4]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_6_io_x_paa = _GEN_59[3]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_6_io_x_eff = _GEN_59[2]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_6_io_x_c = _GEN_59[1]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_7_io_x_ppn = _GEN_63[34:15]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_7_io_x_u = _GEN_63[14]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_7_io_x_ae = _GEN_63[12]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_7_io_x_sw = _GEN_63[11]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_7_io_x_sx = _GEN_63[10]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_7_io_x_sr = _GEN_63[9]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_7_io_x_pw = _GEN_63[8]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_7_io_x_px = _GEN_63[7]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_7_io_x_pr = _GEN_63[6]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_7_io_x_ppp = _GEN_63[5]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_7_io_x_pal = _GEN_63[4]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_7_io_x_paa = _GEN_63[3]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_7_io_x_eff = _GEN_63[2]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_7_io_x_c = _GEN_63[1]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_8_io_x_ppn = superpage_entries_0_data_0[34:15]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_8_io_x_u = superpage_entries_0_data_0[14]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_8_io_x_ae = superpage_entries_0_data_0[12]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_8_io_x_sw = superpage_entries_0_data_0[11]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_8_io_x_sx = superpage_entries_0_data_0[10]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_8_io_x_sr = superpage_entries_0_data_0[9]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_8_io_x_pw = superpage_entries_0_data_0[8]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_8_io_x_px = superpage_entries_0_data_0[7]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_8_io_x_pr = superpage_entries_0_data_0[6]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_8_io_x_ppp = superpage_entries_0_data_0[5]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_8_io_x_pal = superpage_entries_0_data_0[4]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_8_io_x_paa = superpage_entries_0_data_0[3]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_8_io_x_eff = superpage_entries_0_data_0[2]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_8_io_x_c = superpage_entries_0_data_0[1]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_9_io_x_ppn = superpage_entries_1_data_0[34:15]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_9_io_x_u = superpage_entries_1_data_0[14]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_9_io_x_ae = superpage_entries_1_data_0[12]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_9_io_x_sw = superpage_entries_1_data_0[11]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_9_io_x_sx = superpage_entries_1_data_0[10]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_9_io_x_sr = superpage_entries_1_data_0[9]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_9_io_x_pw = superpage_entries_1_data_0[8]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_9_io_x_px = superpage_entries_1_data_0[7]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_9_io_x_pr = superpage_entries_1_data_0[6]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_9_io_x_ppp = superpage_entries_1_data_0[5]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_9_io_x_pal = superpage_entries_1_data_0[4]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_9_io_x_paa = superpage_entries_1_data_0[3]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_9_io_x_eff = superpage_entries_1_data_0[2]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_9_io_x_c = superpage_entries_1_data_0[1]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_10_io_x_ppn = superpage_entries_2_data_0[34:15]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_10_io_x_u = superpage_entries_2_data_0[14]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_10_io_x_ae = superpage_entries_2_data_0[12]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_10_io_x_sw = superpage_entries_2_data_0[11]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_10_io_x_sx = superpage_entries_2_data_0[10]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_10_io_x_sr = superpage_entries_2_data_0[9]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_10_io_x_pw = superpage_entries_2_data_0[8]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_10_io_x_px = superpage_entries_2_data_0[7]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_10_io_x_pr = superpage_entries_2_data_0[6]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_10_io_x_ppp = superpage_entries_2_data_0[5]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_10_io_x_pal = superpage_entries_2_data_0[4]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_10_io_x_paa = superpage_entries_2_data_0[3]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_10_io_x_eff = superpage_entries_2_data_0[2]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_10_io_x_c = superpage_entries_2_data_0[1]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_11_io_x_ppn = superpage_entries_3_data_0[34:15]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_11_io_x_u = superpage_entries_3_data_0[14]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_11_io_x_ae = superpage_entries_3_data_0[12]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_11_io_x_sw = superpage_entries_3_data_0[11]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_11_io_x_sx = superpage_entries_3_data_0[10]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_11_io_x_sr = superpage_entries_3_data_0[9]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_11_io_x_pw = superpage_entries_3_data_0[8]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_11_io_x_px = superpage_entries_3_data_0[7]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_11_io_x_pr = superpage_entries_3_data_0[6]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_11_io_x_ppp = superpage_entries_3_data_0[5]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_11_io_x_pal = superpage_entries_3_data_0[4]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_11_io_x_paa = superpage_entries_3_data_0[3]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_11_io_x_eff = superpage_entries_3_data_0[2]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_11_io_x_c = superpage_entries_3_data_0[1]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_12_io_x_ppn = special_entry_data_0[34:15]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_12_io_x_u = special_entry_data_0[14]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_12_io_x_ae = special_entry_data_0[12]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_12_io_x_sw = special_entry_data_0[11]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_12_io_x_sx = special_entry_data_0[10]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_12_io_x_sr = special_entry_data_0[9]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_12_io_x_pw = special_entry_data_0[8]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_12_io_x_px = special_entry_data_0[7]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_12_io_x_pr = special_entry_data_0[6]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_12_io_x_ppp = special_entry_data_0[5]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_12_io_x_pal = special_entry_data_0[4]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_12_io_x_paa = special_entry_data_0[3]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_12_io_x_eff = special_entry_data_0[2]; // @[TLB.scala 86:77]
  assign ppn_data_barrier_12_io_x_c = special_entry_data_0[1]; // @[TLB.scala 86:77]
  assign entries_barrier_io_x_ppn = _GEN_35[34:15]; // @[TLB.scala 86:77]
  assign entries_barrier_io_x_u = _GEN_35[14]; // @[TLB.scala 86:77]
  assign entries_barrier_io_x_ae = _GEN_35[12]; // @[TLB.scala 86:77]
  assign entries_barrier_io_x_sw = _GEN_35[11]; // @[TLB.scala 86:77]
  assign entries_barrier_io_x_sx = _GEN_35[10]; // @[TLB.scala 86:77]
  assign entries_barrier_io_x_sr = _GEN_35[9]; // @[TLB.scala 86:77]
  assign entries_barrier_io_x_pw = _GEN_35[8]; // @[TLB.scala 86:77]
  assign entries_barrier_io_x_px = _GEN_35[7]; // @[TLB.scala 86:77]
  assign entries_barrier_io_x_pr = _GEN_35[6]; // @[TLB.scala 86:77]
  assign entries_barrier_io_x_ppp = _GEN_35[5]; // @[TLB.scala 86:77]
  assign entries_barrier_io_x_pal = _GEN_35[4]; // @[TLB.scala 86:77]
  assign entries_barrier_io_x_paa = _GEN_35[3]; // @[TLB.scala 86:77]
  assign entries_barrier_io_x_eff = _GEN_35[2]; // @[TLB.scala 86:77]
  assign entries_barrier_io_x_c = _GEN_35[1]; // @[TLB.scala 86:77]
  assign entries_barrier_1_io_x_ppn = _GEN_39[34:15]; // @[TLB.scala 86:77]
  assign entries_barrier_1_io_x_u = _GEN_39[14]; // @[TLB.scala 86:77]
  assign entries_barrier_1_io_x_ae = _GEN_39[12]; // @[TLB.scala 86:77]
  assign entries_barrier_1_io_x_sw = _GEN_39[11]; // @[TLB.scala 86:77]
  assign entries_barrier_1_io_x_sx = _GEN_39[10]; // @[TLB.scala 86:77]
  assign entries_barrier_1_io_x_sr = _GEN_39[9]; // @[TLB.scala 86:77]
  assign entries_barrier_1_io_x_pw = _GEN_39[8]; // @[TLB.scala 86:77]
  assign entries_barrier_1_io_x_px = _GEN_39[7]; // @[TLB.scala 86:77]
  assign entries_barrier_1_io_x_pr = _GEN_39[6]; // @[TLB.scala 86:77]
  assign entries_barrier_1_io_x_ppp = _GEN_39[5]; // @[TLB.scala 86:77]
  assign entries_barrier_1_io_x_pal = _GEN_39[4]; // @[TLB.scala 86:77]
  assign entries_barrier_1_io_x_paa = _GEN_39[3]; // @[TLB.scala 86:77]
  assign entries_barrier_1_io_x_eff = _GEN_39[2]; // @[TLB.scala 86:77]
  assign entries_barrier_1_io_x_c = _GEN_39[1]; // @[TLB.scala 86:77]
  assign entries_barrier_2_io_x_ppn = _GEN_43[34:15]; // @[TLB.scala 86:77]
  assign entries_barrier_2_io_x_u = _GEN_43[14]; // @[TLB.scala 86:77]
  assign entries_barrier_2_io_x_ae = _GEN_43[12]; // @[TLB.scala 86:77]
  assign entries_barrier_2_io_x_sw = _GEN_43[11]; // @[TLB.scala 86:77]
  assign entries_barrier_2_io_x_sx = _GEN_43[10]; // @[TLB.scala 86:77]
  assign entries_barrier_2_io_x_sr = _GEN_43[9]; // @[TLB.scala 86:77]
  assign entries_barrier_2_io_x_pw = _GEN_43[8]; // @[TLB.scala 86:77]
  assign entries_barrier_2_io_x_px = _GEN_43[7]; // @[TLB.scala 86:77]
  assign entries_barrier_2_io_x_pr = _GEN_43[6]; // @[TLB.scala 86:77]
  assign entries_barrier_2_io_x_ppp = _GEN_43[5]; // @[TLB.scala 86:77]
  assign entries_barrier_2_io_x_pal = _GEN_43[4]; // @[TLB.scala 86:77]
  assign entries_barrier_2_io_x_paa = _GEN_43[3]; // @[TLB.scala 86:77]
  assign entries_barrier_2_io_x_eff = _GEN_43[2]; // @[TLB.scala 86:77]
  assign entries_barrier_2_io_x_c = _GEN_43[1]; // @[TLB.scala 86:77]
  assign entries_barrier_3_io_x_ppn = _GEN_47[34:15]; // @[TLB.scala 86:77]
  assign entries_barrier_3_io_x_u = _GEN_47[14]; // @[TLB.scala 86:77]
  assign entries_barrier_3_io_x_ae = _GEN_47[12]; // @[TLB.scala 86:77]
  assign entries_barrier_3_io_x_sw = _GEN_47[11]; // @[TLB.scala 86:77]
  assign entries_barrier_3_io_x_sx = _GEN_47[10]; // @[TLB.scala 86:77]
  assign entries_barrier_3_io_x_sr = _GEN_47[9]; // @[TLB.scala 86:77]
  assign entries_barrier_3_io_x_pw = _GEN_47[8]; // @[TLB.scala 86:77]
  assign entries_barrier_3_io_x_px = _GEN_47[7]; // @[TLB.scala 86:77]
  assign entries_barrier_3_io_x_pr = _GEN_47[6]; // @[TLB.scala 86:77]
  assign entries_barrier_3_io_x_ppp = _GEN_47[5]; // @[TLB.scala 86:77]
  assign entries_barrier_3_io_x_pal = _GEN_47[4]; // @[TLB.scala 86:77]
  assign entries_barrier_3_io_x_paa = _GEN_47[3]; // @[TLB.scala 86:77]
  assign entries_barrier_3_io_x_eff = _GEN_47[2]; // @[TLB.scala 86:77]
  assign entries_barrier_3_io_x_c = _GEN_47[1]; // @[TLB.scala 86:77]
  assign entries_barrier_4_io_x_ppn = _GEN_51[34:15]; // @[TLB.scala 86:77]
  assign entries_barrier_4_io_x_u = _GEN_51[14]; // @[TLB.scala 86:77]
  assign entries_barrier_4_io_x_ae = _GEN_51[12]; // @[TLB.scala 86:77]
  assign entries_barrier_4_io_x_sw = _GEN_51[11]; // @[TLB.scala 86:77]
  assign entries_barrier_4_io_x_sx = _GEN_51[10]; // @[TLB.scala 86:77]
  assign entries_barrier_4_io_x_sr = _GEN_51[9]; // @[TLB.scala 86:77]
  assign entries_barrier_4_io_x_pw = _GEN_51[8]; // @[TLB.scala 86:77]
  assign entries_barrier_4_io_x_px = _GEN_51[7]; // @[TLB.scala 86:77]
  assign entries_barrier_4_io_x_pr = _GEN_51[6]; // @[TLB.scala 86:77]
  assign entries_barrier_4_io_x_ppp = _GEN_51[5]; // @[TLB.scala 86:77]
  assign entries_barrier_4_io_x_pal = _GEN_51[4]; // @[TLB.scala 86:77]
  assign entries_barrier_4_io_x_paa = _GEN_51[3]; // @[TLB.scala 86:77]
  assign entries_barrier_4_io_x_eff = _GEN_51[2]; // @[TLB.scala 86:77]
  assign entries_barrier_4_io_x_c = _GEN_51[1]; // @[TLB.scala 86:77]
  assign entries_barrier_5_io_x_ppn = _GEN_55[34:15]; // @[TLB.scala 86:77]
  assign entries_barrier_5_io_x_u = _GEN_55[14]; // @[TLB.scala 86:77]
  assign entries_barrier_5_io_x_ae = _GEN_55[12]; // @[TLB.scala 86:77]
  assign entries_barrier_5_io_x_sw = _GEN_55[11]; // @[TLB.scala 86:77]
  assign entries_barrier_5_io_x_sx = _GEN_55[10]; // @[TLB.scala 86:77]
  assign entries_barrier_5_io_x_sr = _GEN_55[9]; // @[TLB.scala 86:77]
  assign entries_barrier_5_io_x_pw = _GEN_55[8]; // @[TLB.scala 86:77]
  assign entries_barrier_5_io_x_px = _GEN_55[7]; // @[TLB.scala 86:77]
  assign entries_barrier_5_io_x_pr = _GEN_55[6]; // @[TLB.scala 86:77]
  assign entries_barrier_5_io_x_ppp = _GEN_55[5]; // @[TLB.scala 86:77]
  assign entries_barrier_5_io_x_pal = _GEN_55[4]; // @[TLB.scala 86:77]
  assign entries_barrier_5_io_x_paa = _GEN_55[3]; // @[TLB.scala 86:77]
  assign entries_barrier_5_io_x_eff = _GEN_55[2]; // @[TLB.scala 86:77]
  assign entries_barrier_5_io_x_c = _GEN_55[1]; // @[TLB.scala 86:77]
  assign entries_barrier_6_io_x_ppn = _GEN_59[34:15]; // @[TLB.scala 86:77]
  assign entries_barrier_6_io_x_u = _GEN_59[14]; // @[TLB.scala 86:77]
  assign entries_barrier_6_io_x_ae = _GEN_59[12]; // @[TLB.scala 86:77]
  assign entries_barrier_6_io_x_sw = _GEN_59[11]; // @[TLB.scala 86:77]
  assign entries_barrier_6_io_x_sx = _GEN_59[10]; // @[TLB.scala 86:77]
  assign entries_barrier_6_io_x_sr = _GEN_59[9]; // @[TLB.scala 86:77]
  assign entries_barrier_6_io_x_pw = _GEN_59[8]; // @[TLB.scala 86:77]
  assign entries_barrier_6_io_x_px = _GEN_59[7]; // @[TLB.scala 86:77]
  assign entries_barrier_6_io_x_pr = _GEN_59[6]; // @[TLB.scala 86:77]
  assign entries_barrier_6_io_x_ppp = _GEN_59[5]; // @[TLB.scala 86:77]
  assign entries_barrier_6_io_x_pal = _GEN_59[4]; // @[TLB.scala 86:77]
  assign entries_barrier_6_io_x_paa = _GEN_59[3]; // @[TLB.scala 86:77]
  assign entries_barrier_6_io_x_eff = _GEN_59[2]; // @[TLB.scala 86:77]
  assign entries_barrier_6_io_x_c = _GEN_59[1]; // @[TLB.scala 86:77]
  assign entries_barrier_7_io_x_ppn = _GEN_63[34:15]; // @[TLB.scala 86:77]
  assign entries_barrier_7_io_x_u = _GEN_63[14]; // @[TLB.scala 86:77]
  assign entries_barrier_7_io_x_ae = _GEN_63[12]; // @[TLB.scala 86:77]
  assign entries_barrier_7_io_x_sw = _GEN_63[11]; // @[TLB.scala 86:77]
  assign entries_barrier_7_io_x_sx = _GEN_63[10]; // @[TLB.scala 86:77]
  assign entries_barrier_7_io_x_sr = _GEN_63[9]; // @[TLB.scala 86:77]
  assign entries_barrier_7_io_x_pw = _GEN_63[8]; // @[TLB.scala 86:77]
  assign entries_barrier_7_io_x_px = _GEN_63[7]; // @[TLB.scala 86:77]
  assign entries_barrier_7_io_x_pr = _GEN_63[6]; // @[TLB.scala 86:77]
  assign entries_barrier_7_io_x_ppp = _GEN_63[5]; // @[TLB.scala 86:77]
  assign entries_barrier_7_io_x_pal = _GEN_63[4]; // @[TLB.scala 86:77]
  assign entries_barrier_7_io_x_paa = _GEN_63[3]; // @[TLB.scala 86:77]
  assign entries_barrier_7_io_x_eff = _GEN_63[2]; // @[TLB.scala 86:77]
  assign entries_barrier_7_io_x_c = _GEN_63[1]; // @[TLB.scala 86:77]
  assign entries_barrier_8_io_x_ppn = superpage_entries_0_data_0[34:15]; // @[TLB.scala 86:77]
  assign entries_barrier_8_io_x_u = superpage_entries_0_data_0[14]; // @[TLB.scala 86:77]
  assign entries_barrier_8_io_x_ae = superpage_entries_0_data_0[12]; // @[TLB.scala 86:77]
  assign entries_barrier_8_io_x_sw = superpage_entries_0_data_0[11]; // @[TLB.scala 86:77]
  assign entries_barrier_8_io_x_sx = superpage_entries_0_data_0[10]; // @[TLB.scala 86:77]
  assign entries_barrier_8_io_x_sr = superpage_entries_0_data_0[9]; // @[TLB.scala 86:77]
  assign entries_barrier_8_io_x_pw = superpage_entries_0_data_0[8]; // @[TLB.scala 86:77]
  assign entries_barrier_8_io_x_px = superpage_entries_0_data_0[7]; // @[TLB.scala 86:77]
  assign entries_barrier_8_io_x_pr = superpage_entries_0_data_0[6]; // @[TLB.scala 86:77]
  assign entries_barrier_8_io_x_ppp = superpage_entries_0_data_0[5]; // @[TLB.scala 86:77]
  assign entries_barrier_8_io_x_pal = superpage_entries_0_data_0[4]; // @[TLB.scala 86:77]
  assign entries_barrier_8_io_x_paa = superpage_entries_0_data_0[3]; // @[TLB.scala 86:77]
  assign entries_barrier_8_io_x_eff = superpage_entries_0_data_0[2]; // @[TLB.scala 86:77]
  assign entries_barrier_8_io_x_c = superpage_entries_0_data_0[1]; // @[TLB.scala 86:77]
  assign entries_barrier_9_io_x_ppn = superpage_entries_1_data_0[34:15]; // @[TLB.scala 86:77]
  assign entries_barrier_9_io_x_u = superpage_entries_1_data_0[14]; // @[TLB.scala 86:77]
  assign entries_barrier_9_io_x_ae = superpage_entries_1_data_0[12]; // @[TLB.scala 86:77]
  assign entries_barrier_9_io_x_sw = superpage_entries_1_data_0[11]; // @[TLB.scala 86:77]
  assign entries_barrier_9_io_x_sx = superpage_entries_1_data_0[10]; // @[TLB.scala 86:77]
  assign entries_barrier_9_io_x_sr = superpage_entries_1_data_0[9]; // @[TLB.scala 86:77]
  assign entries_barrier_9_io_x_pw = superpage_entries_1_data_0[8]; // @[TLB.scala 86:77]
  assign entries_barrier_9_io_x_px = superpage_entries_1_data_0[7]; // @[TLB.scala 86:77]
  assign entries_barrier_9_io_x_pr = superpage_entries_1_data_0[6]; // @[TLB.scala 86:77]
  assign entries_barrier_9_io_x_ppp = superpage_entries_1_data_0[5]; // @[TLB.scala 86:77]
  assign entries_barrier_9_io_x_pal = superpage_entries_1_data_0[4]; // @[TLB.scala 86:77]
  assign entries_barrier_9_io_x_paa = superpage_entries_1_data_0[3]; // @[TLB.scala 86:77]
  assign entries_barrier_9_io_x_eff = superpage_entries_1_data_0[2]; // @[TLB.scala 86:77]
  assign entries_barrier_9_io_x_c = superpage_entries_1_data_0[1]; // @[TLB.scala 86:77]
  assign entries_barrier_10_io_x_ppn = superpage_entries_2_data_0[34:15]; // @[TLB.scala 86:77]
  assign entries_barrier_10_io_x_u = superpage_entries_2_data_0[14]; // @[TLB.scala 86:77]
  assign entries_barrier_10_io_x_ae = superpage_entries_2_data_0[12]; // @[TLB.scala 86:77]
  assign entries_barrier_10_io_x_sw = superpage_entries_2_data_0[11]; // @[TLB.scala 86:77]
  assign entries_barrier_10_io_x_sx = superpage_entries_2_data_0[10]; // @[TLB.scala 86:77]
  assign entries_barrier_10_io_x_sr = superpage_entries_2_data_0[9]; // @[TLB.scala 86:77]
  assign entries_barrier_10_io_x_pw = superpage_entries_2_data_0[8]; // @[TLB.scala 86:77]
  assign entries_barrier_10_io_x_px = superpage_entries_2_data_0[7]; // @[TLB.scala 86:77]
  assign entries_barrier_10_io_x_pr = superpage_entries_2_data_0[6]; // @[TLB.scala 86:77]
  assign entries_barrier_10_io_x_ppp = superpage_entries_2_data_0[5]; // @[TLB.scala 86:77]
  assign entries_barrier_10_io_x_pal = superpage_entries_2_data_0[4]; // @[TLB.scala 86:77]
  assign entries_barrier_10_io_x_paa = superpage_entries_2_data_0[3]; // @[TLB.scala 86:77]
  assign entries_barrier_10_io_x_eff = superpage_entries_2_data_0[2]; // @[TLB.scala 86:77]
  assign entries_barrier_10_io_x_c = superpage_entries_2_data_0[1]; // @[TLB.scala 86:77]
  assign entries_barrier_11_io_x_ppn = superpage_entries_3_data_0[34:15]; // @[TLB.scala 86:77]
  assign entries_barrier_11_io_x_u = superpage_entries_3_data_0[14]; // @[TLB.scala 86:77]
  assign entries_barrier_11_io_x_ae = superpage_entries_3_data_0[12]; // @[TLB.scala 86:77]
  assign entries_barrier_11_io_x_sw = superpage_entries_3_data_0[11]; // @[TLB.scala 86:77]
  assign entries_barrier_11_io_x_sx = superpage_entries_3_data_0[10]; // @[TLB.scala 86:77]
  assign entries_barrier_11_io_x_sr = superpage_entries_3_data_0[9]; // @[TLB.scala 86:77]
  assign entries_barrier_11_io_x_pw = superpage_entries_3_data_0[8]; // @[TLB.scala 86:77]
  assign entries_barrier_11_io_x_px = superpage_entries_3_data_0[7]; // @[TLB.scala 86:77]
  assign entries_barrier_11_io_x_pr = superpage_entries_3_data_0[6]; // @[TLB.scala 86:77]
  assign entries_barrier_11_io_x_ppp = superpage_entries_3_data_0[5]; // @[TLB.scala 86:77]
  assign entries_barrier_11_io_x_pal = superpage_entries_3_data_0[4]; // @[TLB.scala 86:77]
  assign entries_barrier_11_io_x_paa = superpage_entries_3_data_0[3]; // @[TLB.scala 86:77]
  assign entries_barrier_11_io_x_eff = superpage_entries_3_data_0[2]; // @[TLB.scala 86:77]
  assign entries_barrier_11_io_x_c = superpage_entries_3_data_0[1]; // @[TLB.scala 86:77]
  assign entries_barrier_12_io_x_ppn = special_entry_data_0[34:15]; // @[TLB.scala 86:77]
  assign entries_barrier_12_io_x_u = special_entry_data_0[14]; // @[TLB.scala 86:77]
  assign entries_barrier_12_io_x_ae = special_entry_data_0[12]; // @[TLB.scala 86:77]
  assign entries_barrier_12_io_x_sw = special_entry_data_0[11]; // @[TLB.scala 86:77]
  assign entries_barrier_12_io_x_sx = special_entry_data_0[10]; // @[TLB.scala 86:77]
  assign entries_barrier_12_io_x_sr = special_entry_data_0[9]; // @[TLB.scala 86:77]
  assign entries_barrier_12_io_x_pw = special_entry_data_0[8]; // @[TLB.scala 86:77]
  assign entries_barrier_12_io_x_px = special_entry_data_0[7]; // @[TLB.scala 86:77]
  assign entries_barrier_12_io_x_pr = special_entry_data_0[6]; // @[TLB.scala 86:77]
  assign entries_barrier_12_io_x_ppp = special_entry_data_0[5]; // @[TLB.scala 86:77]
  assign entries_barrier_12_io_x_pal = special_entry_data_0[4]; // @[TLB.scala 86:77]
  assign entries_barrier_12_io_x_paa = special_entry_data_0[3]; // @[TLB.scala 86:77]
  assign entries_barrier_12_io_x_eff = special_entry_data_0[2]; // @[TLB.scala 86:77]
  assign entries_barrier_12_io_x_c = special_entry_data_0[1]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_io_x_ppn = _GEN_35[34:15]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_io_x_u = _GEN_35[14]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_io_x_ae = _GEN_35[12]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_io_x_sw = _GEN_35[11]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_io_x_sx = _GEN_35[10]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_io_x_sr = _GEN_35[9]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_io_x_pw = _GEN_35[8]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_io_x_px = _GEN_35[7]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_io_x_pr = _GEN_35[6]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_io_x_ppp = _GEN_35[5]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_io_x_pal = _GEN_35[4]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_io_x_paa = _GEN_35[3]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_io_x_eff = _GEN_35[2]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_io_x_c = _GEN_35[1]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_1_io_x_ppn = _GEN_39[34:15]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_1_io_x_u = _GEN_39[14]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_1_io_x_ae = _GEN_39[12]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_1_io_x_sw = _GEN_39[11]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_1_io_x_sx = _GEN_39[10]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_1_io_x_sr = _GEN_39[9]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_1_io_x_pw = _GEN_39[8]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_1_io_x_px = _GEN_39[7]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_1_io_x_pr = _GEN_39[6]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_1_io_x_ppp = _GEN_39[5]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_1_io_x_pal = _GEN_39[4]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_1_io_x_paa = _GEN_39[3]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_1_io_x_eff = _GEN_39[2]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_1_io_x_c = _GEN_39[1]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_2_io_x_ppn = _GEN_43[34:15]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_2_io_x_u = _GEN_43[14]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_2_io_x_ae = _GEN_43[12]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_2_io_x_sw = _GEN_43[11]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_2_io_x_sx = _GEN_43[10]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_2_io_x_sr = _GEN_43[9]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_2_io_x_pw = _GEN_43[8]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_2_io_x_px = _GEN_43[7]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_2_io_x_pr = _GEN_43[6]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_2_io_x_ppp = _GEN_43[5]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_2_io_x_pal = _GEN_43[4]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_2_io_x_paa = _GEN_43[3]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_2_io_x_eff = _GEN_43[2]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_2_io_x_c = _GEN_43[1]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_3_io_x_ppn = _GEN_47[34:15]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_3_io_x_u = _GEN_47[14]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_3_io_x_ae = _GEN_47[12]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_3_io_x_sw = _GEN_47[11]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_3_io_x_sx = _GEN_47[10]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_3_io_x_sr = _GEN_47[9]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_3_io_x_pw = _GEN_47[8]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_3_io_x_px = _GEN_47[7]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_3_io_x_pr = _GEN_47[6]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_3_io_x_ppp = _GEN_47[5]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_3_io_x_pal = _GEN_47[4]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_3_io_x_paa = _GEN_47[3]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_3_io_x_eff = _GEN_47[2]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_3_io_x_c = _GEN_47[1]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_4_io_x_ppn = _GEN_51[34:15]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_4_io_x_u = _GEN_51[14]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_4_io_x_ae = _GEN_51[12]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_4_io_x_sw = _GEN_51[11]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_4_io_x_sx = _GEN_51[10]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_4_io_x_sr = _GEN_51[9]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_4_io_x_pw = _GEN_51[8]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_4_io_x_px = _GEN_51[7]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_4_io_x_pr = _GEN_51[6]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_4_io_x_ppp = _GEN_51[5]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_4_io_x_pal = _GEN_51[4]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_4_io_x_paa = _GEN_51[3]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_4_io_x_eff = _GEN_51[2]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_4_io_x_c = _GEN_51[1]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_5_io_x_ppn = _GEN_55[34:15]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_5_io_x_u = _GEN_55[14]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_5_io_x_ae = _GEN_55[12]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_5_io_x_sw = _GEN_55[11]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_5_io_x_sx = _GEN_55[10]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_5_io_x_sr = _GEN_55[9]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_5_io_x_pw = _GEN_55[8]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_5_io_x_px = _GEN_55[7]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_5_io_x_pr = _GEN_55[6]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_5_io_x_ppp = _GEN_55[5]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_5_io_x_pal = _GEN_55[4]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_5_io_x_paa = _GEN_55[3]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_5_io_x_eff = _GEN_55[2]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_5_io_x_c = _GEN_55[1]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_6_io_x_ppn = _GEN_59[34:15]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_6_io_x_u = _GEN_59[14]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_6_io_x_ae = _GEN_59[12]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_6_io_x_sw = _GEN_59[11]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_6_io_x_sx = _GEN_59[10]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_6_io_x_sr = _GEN_59[9]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_6_io_x_pw = _GEN_59[8]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_6_io_x_px = _GEN_59[7]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_6_io_x_pr = _GEN_59[6]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_6_io_x_ppp = _GEN_59[5]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_6_io_x_pal = _GEN_59[4]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_6_io_x_paa = _GEN_59[3]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_6_io_x_eff = _GEN_59[2]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_6_io_x_c = _GEN_59[1]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_7_io_x_ppn = _GEN_63[34:15]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_7_io_x_u = _GEN_63[14]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_7_io_x_ae = _GEN_63[12]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_7_io_x_sw = _GEN_63[11]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_7_io_x_sx = _GEN_63[10]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_7_io_x_sr = _GEN_63[9]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_7_io_x_pw = _GEN_63[8]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_7_io_x_px = _GEN_63[7]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_7_io_x_pr = _GEN_63[6]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_7_io_x_ppp = _GEN_63[5]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_7_io_x_pal = _GEN_63[4]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_7_io_x_paa = _GEN_63[3]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_7_io_x_eff = _GEN_63[2]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_7_io_x_c = _GEN_63[1]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_8_io_x_ppn = superpage_entries_0_data_0[34:15]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_8_io_x_u = superpage_entries_0_data_0[14]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_8_io_x_ae = superpage_entries_0_data_0[12]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_8_io_x_sw = superpage_entries_0_data_0[11]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_8_io_x_sx = superpage_entries_0_data_0[10]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_8_io_x_sr = superpage_entries_0_data_0[9]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_8_io_x_pw = superpage_entries_0_data_0[8]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_8_io_x_px = superpage_entries_0_data_0[7]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_8_io_x_pr = superpage_entries_0_data_0[6]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_8_io_x_ppp = superpage_entries_0_data_0[5]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_8_io_x_pal = superpage_entries_0_data_0[4]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_8_io_x_paa = superpage_entries_0_data_0[3]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_8_io_x_eff = superpage_entries_0_data_0[2]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_8_io_x_c = superpage_entries_0_data_0[1]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_9_io_x_ppn = superpage_entries_1_data_0[34:15]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_9_io_x_u = superpage_entries_1_data_0[14]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_9_io_x_ae = superpage_entries_1_data_0[12]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_9_io_x_sw = superpage_entries_1_data_0[11]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_9_io_x_sx = superpage_entries_1_data_0[10]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_9_io_x_sr = superpage_entries_1_data_0[9]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_9_io_x_pw = superpage_entries_1_data_0[8]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_9_io_x_px = superpage_entries_1_data_0[7]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_9_io_x_pr = superpage_entries_1_data_0[6]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_9_io_x_ppp = superpage_entries_1_data_0[5]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_9_io_x_pal = superpage_entries_1_data_0[4]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_9_io_x_paa = superpage_entries_1_data_0[3]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_9_io_x_eff = superpage_entries_1_data_0[2]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_9_io_x_c = superpage_entries_1_data_0[1]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_10_io_x_ppn = superpage_entries_2_data_0[34:15]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_10_io_x_u = superpage_entries_2_data_0[14]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_10_io_x_ae = superpage_entries_2_data_0[12]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_10_io_x_sw = superpage_entries_2_data_0[11]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_10_io_x_sx = superpage_entries_2_data_0[10]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_10_io_x_sr = superpage_entries_2_data_0[9]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_10_io_x_pw = superpage_entries_2_data_0[8]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_10_io_x_px = superpage_entries_2_data_0[7]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_10_io_x_pr = superpage_entries_2_data_0[6]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_10_io_x_ppp = superpage_entries_2_data_0[5]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_10_io_x_pal = superpage_entries_2_data_0[4]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_10_io_x_paa = superpage_entries_2_data_0[3]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_10_io_x_eff = superpage_entries_2_data_0[2]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_10_io_x_c = superpage_entries_2_data_0[1]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_11_io_x_ppn = superpage_entries_3_data_0[34:15]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_11_io_x_u = superpage_entries_3_data_0[14]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_11_io_x_ae = superpage_entries_3_data_0[12]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_11_io_x_sw = superpage_entries_3_data_0[11]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_11_io_x_sx = superpage_entries_3_data_0[10]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_11_io_x_sr = superpage_entries_3_data_0[9]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_11_io_x_pw = superpage_entries_3_data_0[8]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_11_io_x_px = superpage_entries_3_data_0[7]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_11_io_x_pr = superpage_entries_3_data_0[6]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_11_io_x_ppp = superpage_entries_3_data_0[5]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_11_io_x_pal = superpage_entries_3_data_0[4]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_11_io_x_paa = superpage_entries_3_data_0[3]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_11_io_x_eff = superpage_entries_3_data_0[2]; // @[TLB.scala 86:77]
  assign normal_entries_barrier_11_io_x_c = superpage_entries_3_data_0[1]; // @[TLB.scala 86:77]
  always @(posedge clock) begin
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_7) begin // @[TLB.scala 249:72]
            sectored_entries_0_tag <= r_refill_tag; // @[TLB.scala 118:14]
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_7) begin // @[TLB.scala 249:72]
            sectored_entries_0_data_0 <= _GEN_89;
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_7) begin // @[TLB.scala 249:72]
            sectored_entries_0_data_1 <= _GEN_90;
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_7) begin // @[TLB.scala 249:72]
            sectored_entries_0_data_2 <= _GEN_91;
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_7) begin // @[TLB.scala 249:72]
            sectored_entries_0_data_3 <= _GEN_92;
          end
        end
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      sectored_entries_0_valid_0 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (_T_59) begin // @[TLB.scala 135:68]
          sectored_entries_0_valid_0 <= _GEN_673;
        end else begin
          sectored_entries_0_valid_0 <= _GEN_669;
        end
      end else begin
        sectored_entries_0_valid_0 <= _GEN_685;
      end
    end else if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        sectored_entries_0_valid_0 <= _GEN_305;
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      sectored_entries_0_valid_1 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (_T_59) begin // @[TLB.scala 135:68]
          sectored_entries_0_valid_1 <= _GEN_674;
        end else begin
          sectored_entries_0_valid_1 <= _GEN_670;
        end
      end else begin
        sectored_entries_0_valid_1 <= _GEN_686;
      end
    end else if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        sectored_entries_0_valid_1 <= _GEN_306;
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      sectored_entries_0_valid_2 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (_T_59) begin // @[TLB.scala 135:68]
          sectored_entries_0_valid_2 <= _GEN_675;
        end else begin
          sectored_entries_0_valid_2 <= _GEN_671;
        end
      end else begin
        sectored_entries_0_valid_2 <= _GEN_687;
      end
    end else if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        sectored_entries_0_valid_2 <= _GEN_307;
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      sectored_entries_0_valid_3 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (_T_59) begin // @[TLB.scala 135:68]
          sectored_entries_0_valid_3 <= _GEN_676;
        end else begin
          sectored_entries_0_valid_3 <= _GEN_672;
        end
      end else begin
        sectored_entries_0_valid_3 <= _GEN_688;
      end
    end else if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        sectored_entries_0_valid_3 <= _GEN_308;
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_9) begin // @[TLB.scala 249:72]
            sectored_entries_1_tag <= r_refill_tag; // @[TLB.scala 118:14]
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_9) begin // @[TLB.scala 249:72]
            sectored_entries_1_data_0 <= _GEN_115;
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_9) begin // @[TLB.scala 249:72]
            sectored_entries_1_data_1 <= _GEN_116;
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_9) begin // @[TLB.scala 249:72]
            sectored_entries_1_data_2 <= _GEN_117;
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_9) begin // @[TLB.scala 249:72]
            sectored_entries_1_data_3 <= _GEN_118;
          end
        end
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      sectored_entries_1_valid_0 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (_T_198) begin // @[TLB.scala 135:68]
          sectored_entries_1_valid_0 <= _GEN_701;
        end else begin
          sectored_entries_1_valid_0 <= _GEN_697;
        end
      end else begin
        sectored_entries_1_valid_0 <= _GEN_713;
      end
    end else if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        sectored_entries_1_valid_0 <= _GEN_315;
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      sectored_entries_1_valid_1 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (_T_198) begin // @[TLB.scala 135:68]
          sectored_entries_1_valid_1 <= _GEN_702;
        end else begin
          sectored_entries_1_valid_1 <= _GEN_698;
        end
      end else begin
        sectored_entries_1_valid_1 <= _GEN_714;
      end
    end else if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        sectored_entries_1_valid_1 <= _GEN_316;
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      sectored_entries_1_valid_2 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (_T_198) begin // @[TLB.scala 135:68]
          sectored_entries_1_valid_2 <= _GEN_703;
        end else begin
          sectored_entries_1_valid_2 <= _GEN_699;
        end
      end else begin
        sectored_entries_1_valid_2 <= _GEN_715;
      end
    end else if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        sectored_entries_1_valid_2 <= _GEN_317;
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      sectored_entries_1_valid_3 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (_T_198) begin // @[TLB.scala 135:68]
          sectored_entries_1_valid_3 <= _GEN_704;
        end else begin
          sectored_entries_1_valid_3 <= _GEN_700;
        end
      end else begin
        sectored_entries_1_valid_3 <= _GEN_716;
      end
    end else if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        sectored_entries_1_valid_3 <= _GEN_318;
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_11) begin // @[TLB.scala 249:72]
            sectored_entries_2_tag <= r_refill_tag; // @[TLB.scala 118:14]
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_11) begin // @[TLB.scala 249:72]
            sectored_entries_2_data_0 <= _GEN_141;
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_11) begin // @[TLB.scala 249:72]
            sectored_entries_2_data_1 <= _GEN_142;
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_11) begin // @[TLB.scala 249:72]
            sectored_entries_2_data_2 <= _GEN_143;
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_11) begin // @[TLB.scala 249:72]
            sectored_entries_2_data_3 <= _GEN_144;
          end
        end
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      sectored_entries_2_valid_0 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (_T_337) begin // @[TLB.scala 135:68]
          sectored_entries_2_valid_0 <= _GEN_729;
        end else begin
          sectored_entries_2_valid_0 <= _GEN_725;
        end
      end else begin
        sectored_entries_2_valid_0 <= _GEN_741;
      end
    end else if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        sectored_entries_2_valid_0 <= _GEN_325;
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      sectored_entries_2_valid_1 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (_T_337) begin // @[TLB.scala 135:68]
          sectored_entries_2_valid_1 <= _GEN_730;
        end else begin
          sectored_entries_2_valid_1 <= _GEN_726;
        end
      end else begin
        sectored_entries_2_valid_1 <= _GEN_742;
      end
    end else if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        sectored_entries_2_valid_1 <= _GEN_326;
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      sectored_entries_2_valid_2 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (_T_337) begin // @[TLB.scala 135:68]
          sectored_entries_2_valid_2 <= _GEN_731;
        end else begin
          sectored_entries_2_valid_2 <= _GEN_727;
        end
      end else begin
        sectored_entries_2_valid_2 <= _GEN_743;
      end
    end else if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        sectored_entries_2_valid_2 <= _GEN_327;
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      sectored_entries_2_valid_3 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (_T_337) begin // @[TLB.scala 135:68]
          sectored_entries_2_valid_3 <= _GEN_732;
        end else begin
          sectored_entries_2_valid_3 <= _GEN_728;
        end
      end else begin
        sectored_entries_2_valid_3 <= _GEN_744;
      end
    end else if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        sectored_entries_2_valid_3 <= _GEN_328;
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_13) begin // @[TLB.scala 249:72]
            sectored_entries_3_tag <= r_refill_tag; // @[TLB.scala 118:14]
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_13) begin // @[TLB.scala 249:72]
            sectored_entries_3_data_0 <= _GEN_167;
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_13) begin // @[TLB.scala 249:72]
            sectored_entries_3_data_1 <= _GEN_168;
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_13) begin // @[TLB.scala 249:72]
            sectored_entries_3_data_2 <= _GEN_169;
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_13) begin // @[TLB.scala 249:72]
            sectored_entries_3_data_3 <= _GEN_170;
          end
        end
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      sectored_entries_3_valid_0 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (_T_476) begin // @[TLB.scala 135:68]
          sectored_entries_3_valid_0 <= _GEN_757;
        end else begin
          sectored_entries_3_valid_0 <= _GEN_753;
        end
      end else begin
        sectored_entries_3_valid_0 <= _GEN_769;
      end
    end else if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        sectored_entries_3_valid_0 <= _GEN_335;
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      sectored_entries_3_valid_1 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (_T_476) begin // @[TLB.scala 135:68]
          sectored_entries_3_valid_1 <= _GEN_758;
        end else begin
          sectored_entries_3_valid_1 <= _GEN_754;
        end
      end else begin
        sectored_entries_3_valid_1 <= _GEN_770;
      end
    end else if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        sectored_entries_3_valid_1 <= _GEN_336;
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      sectored_entries_3_valid_2 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (_T_476) begin // @[TLB.scala 135:68]
          sectored_entries_3_valid_2 <= _GEN_759;
        end else begin
          sectored_entries_3_valid_2 <= _GEN_755;
        end
      end else begin
        sectored_entries_3_valid_2 <= _GEN_771;
      end
    end else if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        sectored_entries_3_valid_2 <= _GEN_337;
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      sectored_entries_3_valid_3 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (_T_476) begin // @[TLB.scala 135:68]
          sectored_entries_3_valid_3 <= _GEN_760;
        end else begin
          sectored_entries_3_valid_3 <= _GEN_756;
        end
      end else begin
        sectored_entries_3_valid_3 <= _GEN_772;
      end
    end else if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        sectored_entries_3_valid_3 <= _GEN_338;
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_15) begin // @[TLB.scala 249:72]
            sectored_entries_4_tag <= r_refill_tag; // @[TLB.scala 118:14]
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_15) begin // @[TLB.scala 249:72]
            sectored_entries_4_data_0 <= _GEN_193;
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_15) begin // @[TLB.scala 249:72]
            sectored_entries_4_data_1 <= _GEN_194;
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_15) begin // @[TLB.scala 249:72]
            sectored_entries_4_data_2 <= _GEN_195;
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_15) begin // @[TLB.scala 249:72]
            sectored_entries_4_data_3 <= _GEN_196;
          end
        end
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      sectored_entries_4_valid_0 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (_T_615) begin // @[TLB.scala 135:68]
          sectored_entries_4_valid_0 <= _GEN_785;
        end else begin
          sectored_entries_4_valid_0 <= _GEN_781;
        end
      end else begin
        sectored_entries_4_valid_0 <= _GEN_797;
      end
    end else if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        sectored_entries_4_valid_0 <= _GEN_345;
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      sectored_entries_4_valid_1 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (_T_615) begin // @[TLB.scala 135:68]
          sectored_entries_4_valid_1 <= _GEN_786;
        end else begin
          sectored_entries_4_valid_1 <= _GEN_782;
        end
      end else begin
        sectored_entries_4_valid_1 <= _GEN_798;
      end
    end else if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        sectored_entries_4_valid_1 <= _GEN_346;
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      sectored_entries_4_valid_2 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (_T_615) begin // @[TLB.scala 135:68]
          sectored_entries_4_valid_2 <= _GEN_787;
        end else begin
          sectored_entries_4_valid_2 <= _GEN_783;
        end
      end else begin
        sectored_entries_4_valid_2 <= _GEN_799;
      end
    end else if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        sectored_entries_4_valid_2 <= _GEN_347;
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      sectored_entries_4_valid_3 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (_T_615) begin // @[TLB.scala 135:68]
          sectored_entries_4_valid_3 <= _GEN_788;
        end else begin
          sectored_entries_4_valid_3 <= _GEN_784;
        end
      end else begin
        sectored_entries_4_valid_3 <= _GEN_800;
      end
    end else if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        sectored_entries_4_valid_3 <= _GEN_348;
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_17) begin // @[TLB.scala 249:72]
            sectored_entries_5_tag <= r_refill_tag; // @[TLB.scala 118:14]
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_17) begin // @[TLB.scala 249:72]
            sectored_entries_5_data_0 <= _GEN_219;
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_17) begin // @[TLB.scala 249:72]
            sectored_entries_5_data_1 <= _GEN_220;
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_17) begin // @[TLB.scala 249:72]
            sectored_entries_5_data_2 <= _GEN_221;
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_17) begin // @[TLB.scala 249:72]
            sectored_entries_5_data_3 <= _GEN_222;
          end
        end
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      sectored_entries_5_valid_0 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (_T_754) begin // @[TLB.scala 135:68]
          sectored_entries_5_valid_0 <= _GEN_813;
        end else begin
          sectored_entries_5_valid_0 <= _GEN_809;
        end
      end else begin
        sectored_entries_5_valid_0 <= _GEN_825;
      end
    end else if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        sectored_entries_5_valid_0 <= _GEN_355;
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      sectored_entries_5_valid_1 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (_T_754) begin // @[TLB.scala 135:68]
          sectored_entries_5_valid_1 <= _GEN_814;
        end else begin
          sectored_entries_5_valid_1 <= _GEN_810;
        end
      end else begin
        sectored_entries_5_valid_1 <= _GEN_826;
      end
    end else if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        sectored_entries_5_valid_1 <= _GEN_356;
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      sectored_entries_5_valid_2 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (_T_754) begin // @[TLB.scala 135:68]
          sectored_entries_5_valid_2 <= _GEN_815;
        end else begin
          sectored_entries_5_valid_2 <= _GEN_811;
        end
      end else begin
        sectored_entries_5_valid_2 <= _GEN_827;
      end
    end else if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        sectored_entries_5_valid_2 <= _GEN_357;
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      sectored_entries_5_valid_3 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (_T_754) begin // @[TLB.scala 135:68]
          sectored_entries_5_valid_3 <= _GEN_816;
        end else begin
          sectored_entries_5_valid_3 <= _GEN_812;
        end
      end else begin
        sectored_entries_5_valid_3 <= _GEN_828;
      end
    end else if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        sectored_entries_5_valid_3 <= _GEN_358;
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_19) begin // @[TLB.scala 249:72]
            sectored_entries_6_tag <= r_refill_tag; // @[TLB.scala 118:14]
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_19) begin // @[TLB.scala 249:72]
            sectored_entries_6_data_0 <= _GEN_245;
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_19) begin // @[TLB.scala 249:72]
            sectored_entries_6_data_1 <= _GEN_246;
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_19) begin // @[TLB.scala 249:72]
            sectored_entries_6_data_2 <= _GEN_247;
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_19) begin // @[TLB.scala 249:72]
            sectored_entries_6_data_3 <= _GEN_248;
          end
        end
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      sectored_entries_6_valid_0 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (_T_893) begin // @[TLB.scala 135:68]
          sectored_entries_6_valid_0 <= _GEN_841;
        end else begin
          sectored_entries_6_valid_0 <= _GEN_837;
        end
      end else begin
        sectored_entries_6_valid_0 <= _GEN_853;
      end
    end else if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        sectored_entries_6_valid_0 <= _GEN_365;
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      sectored_entries_6_valid_1 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (_T_893) begin // @[TLB.scala 135:68]
          sectored_entries_6_valid_1 <= _GEN_842;
        end else begin
          sectored_entries_6_valid_1 <= _GEN_838;
        end
      end else begin
        sectored_entries_6_valid_1 <= _GEN_854;
      end
    end else if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        sectored_entries_6_valid_1 <= _GEN_366;
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      sectored_entries_6_valid_2 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (_T_893) begin // @[TLB.scala 135:68]
          sectored_entries_6_valid_2 <= _GEN_843;
        end else begin
          sectored_entries_6_valid_2 <= _GEN_839;
        end
      end else begin
        sectored_entries_6_valid_2 <= _GEN_855;
      end
    end else if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        sectored_entries_6_valid_2 <= _GEN_367;
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      sectored_entries_6_valid_3 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (_T_893) begin // @[TLB.scala 135:68]
          sectored_entries_6_valid_3 <= _GEN_844;
        end else begin
          sectored_entries_6_valid_3 <= _GEN_840;
        end
      end else begin
        sectored_entries_6_valid_3 <= _GEN_856;
      end
    end else if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        sectored_entries_6_valid_3 <= _GEN_368;
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_21) begin // @[TLB.scala 249:72]
            sectored_entries_7_tag <= r_refill_tag; // @[TLB.scala 118:14]
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_21) begin // @[TLB.scala 249:72]
            sectored_entries_7_data_0 <= _GEN_271;
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_21) begin // @[TLB.scala 249:72]
            sectored_entries_7_data_1 <= _GEN_272;
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_21) begin // @[TLB.scala 249:72]
            sectored_entries_7_data_2 <= _GEN_273;
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (!(_T_2)) begin // @[TLB.scala 242:54]
          if (_T_21) begin // @[TLB.scala 249:72]
            sectored_entries_7_data_3 <= _GEN_274;
          end
        end
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      sectored_entries_7_valid_0 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (_T_1032) begin // @[TLB.scala 135:68]
          sectored_entries_7_valid_0 <= _GEN_869;
        end else begin
          sectored_entries_7_valid_0 <= _GEN_865;
        end
      end else begin
        sectored_entries_7_valid_0 <= _GEN_881;
      end
    end else if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        sectored_entries_7_valid_0 <= _GEN_375;
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      sectored_entries_7_valid_1 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (_T_1032) begin // @[TLB.scala 135:68]
          sectored_entries_7_valid_1 <= _GEN_870;
        end else begin
          sectored_entries_7_valid_1 <= _GEN_866;
        end
      end else begin
        sectored_entries_7_valid_1 <= _GEN_882;
      end
    end else if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        sectored_entries_7_valid_1 <= _GEN_376;
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      sectored_entries_7_valid_2 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (_T_1032) begin // @[TLB.scala 135:68]
          sectored_entries_7_valid_2 <= _GEN_871;
        end else begin
          sectored_entries_7_valid_2 <= _GEN_867;
        end
      end else begin
        sectored_entries_7_valid_2 <= _GEN_883;
      end
    end else if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        sectored_entries_7_valid_2 <= _GEN_377;
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      sectored_entries_7_valid_3 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (_T_1032) begin // @[TLB.scala 135:68]
          sectored_entries_7_valid_3 <= _GEN_872;
        end else begin
          sectored_entries_7_valid_3 <= _GEN_868;
        end
      end else begin
        sectored_entries_7_valid_3 <= _GEN_884;
      end
    end else if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        sectored_entries_7_valid_3 <= _GEN_378;
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (_T_2) begin // @[TLB.scala 242:54]
          if (_T_3) begin // @[TLB.scala 243:89]
            superpage_entries_0_level <= {{1'd0}, io_ptw_resp_bits_level[0]}; // @[TLB.scala 119:16]
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (_T_2) begin // @[TLB.scala 242:54]
          if (_T_3) begin // @[TLB.scala 243:89]
            superpage_entries_0_tag <= r_refill_tag; // @[TLB.scala 118:14]
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (_T_2) begin // @[TLB.scala 242:54]
          if (_T_3) begin // @[TLB.scala 243:89]
            superpage_entries_0_data_0 <= _special_entry_data_0_T; // @[TLB.scala 123:15]
          end
        end
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      superpage_entries_0_valid_0 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (superpage_hits_0) begin // @[TLB.scala 129:23]
          superpage_entries_0_valid_0 <= 1'h0; // @[TLB.scala 126:38]
        end else begin
          superpage_entries_0_valid_0 <= _GEN_491;
        end
      end else begin
        superpage_entries_0_valid_0 <= _GEN_891;
      end
    end else begin
      superpage_entries_0_valid_0 <= _GEN_491;
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (_T_2) begin // @[TLB.scala 242:54]
          if (_T_4) begin // @[TLB.scala 243:89]
            superpage_entries_1_level <= {{1'd0}, io_ptw_resp_bits_level[0]}; // @[TLB.scala 119:16]
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (_T_2) begin // @[TLB.scala 242:54]
          if (_T_4) begin // @[TLB.scala 243:89]
            superpage_entries_1_tag <= r_refill_tag; // @[TLB.scala 118:14]
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (_T_2) begin // @[TLB.scala 242:54]
          if (_T_4) begin // @[TLB.scala 243:89]
            superpage_entries_1_data_0 <= _special_entry_data_0_T; // @[TLB.scala 123:15]
          end
        end
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      superpage_entries_1_valid_0 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (superpage_hits_1) begin // @[TLB.scala 129:23]
          superpage_entries_1_valid_0 <= 1'h0; // @[TLB.scala 126:38]
        end else begin
          superpage_entries_1_valid_0 <= _GEN_495;
        end
      end else begin
        superpage_entries_1_valid_0 <= _GEN_895;
      end
    end else begin
      superpage_entries_1_valid_0 <= _GEN_495;
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (_T_2) begin // @[TLB.scala 242:54]
          if (_T_5) begin // @[TLB.scala 243:89]
            superpage_entries_2_level <= {{1'd0}, io_ptw_resp_bits_level[0]}; // @[TLB.scala 119:16]
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (_T_2) begin // @[TLB.scala 242:54]
          if (_T_5) begin // @[TLB.scala 243:89]
            superpage_entries_2_tag <= r_refill_tag; // @[TLB.scala 118:14]
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (_T_2) begin // @[TLB.scala 242:54]
          if (_T_5) begin // @[TLB.scala 243:89]
            superpage_entries_2_data_0 <= _special_entry_data_0_T; // @[TLB.scala 123:15]
          end
        end
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      superpage_entries_2_valid_0 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (superpage_hits_2) begin // @[TLB.scala 129:23]
          superpage_entries_2_valid_0 <= 1'h0; // @[TLB.scala 126:38]
        end else begin
          superpage_entries_2_valid_0 <= _GEN_499;
        end
      end else begin
        superpage_entries_2_valid_0 <= _GEN_899;
      end
    end else begin
      superpage_entries_2_valid_0 <= _GEN_499;
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (_T_2) begin // @[TLB.scala 242:54]
          if (_T_6) begin // @[TLB.scala 243:89]
            superpage_entries_3_level <= {{1'd0}, io_ptw_resp_bits_level[0]}; // @[TLB.scala 119:16]
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (_T_2) begin // @[TLB.scala 242:54]
          if (_T_6) begin // @[TLB.scala 243:89]
            superpage_entries_3_tag <= r_refill_tag; // @[TLB.scala 118:14]
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (!(_T)) begin // @[TLB.scala 237:68]
        if (_T_2) begin // @[TLB.scala 242:54]
          if (_T_6) begin // @[TLB.scala 243:89]
            superpage_entries_3_data_0 <= _special_entry_data_0_T; // @[TLB.scala 123:15]
          end
        end
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      superpage_entries_3_valid_0 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (superpage_hits_3) begin // @[TLB.scala 129:23]
          superpage_entries_3_valid_0 <= 1'h0; // @[TLB.scala 126:38]
        end else begin
          superpage_entries_3_valid_0 <= _GEN_503;
        end
      end else begin
        superpage_entries_3_valid_0 <= _GEN_903;
      end
    end else begin
      superpage_entries_3_valid_0 <= _GEN_503;
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (_T) begin // @[TLB.scala 237:68]
        special_entry_level <= io_ptw_resp_bits_level; // @[TLB.scala 119:16]
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (_T) begin // @[TLB.scala 237:68]
        special_entry_tag <= r_refill_tag; // @[TLB.scala 118:14]
      end
    end
    if (io_ptw_resp_valid) begin // @[TLB.scala 217:20]
      if (_T) begin // @[TLB.scala 237:68]
        special_entry_data_0 <= _special_entry_data_0_T; // @[TLB.scala 123:15]
      end
    end
    if (_T_1326) begin // @[TLB.scala 388:34]
      special_entry_valid_0 <= 1'h0; // @[TLB.scala 126:38]
    end else if (io_sfence_valid) begin // @[TLB.scala 380:19]
      if (io_sfence_bits_rs1) begin // @[TLB.scala 383:35]
        if (_hitsVec_T_106) begin // @[TLB.scala 129:23]
          special_entry_valid_0 <= 1'h0; // @[TLB.scala 126:38]
        end else begin
          special_entry_valid_0 <= _GEN_487;
        end
      end else begin
        special_entry_valid_0 <= _GEN_907;
      end
    end else begin
      special_entry_valid_0 <= _GEN_487;
    end
    if (reset) begin // @[TLB.scala 169:18]
      state <= 2'h0; // @[TLB.scala 169:18]
    end else if (io_ptw_resp_valid) begin // @[TLB.scala 376:30]
      state <= 2'h0; // @[TLB.scala 377:13]
    end else if (_T_45) begin // @[TLB.scala 373:39]
      state <= 2'h3; // @[TLB.scala 374:13]
    end else if (_invalidate_refill_T) begin // @[TLB.scala 368:32]
      state <= _GEN_661;
    end else begin
      state <= _GEN_653;
    end
    if (_T_42) begin // @[TLB.scala 359:38]
      r_refill_tag <= vpn; // @[TLB.scala 361:20]
    end
    if (_T_42) begin // @[TLB.scala 359:38]
      if (&r_superpage_repl_addr_valids) begin // @[TLB.scala 407:8]
        r_superpage_repl_addr <= _r_superpage_repl_addr_T_2;
      end else if (_r_superpage_repl_addr_T_4[0]) begin // @[Mux.scala 47:69]
        r_superpage_repl_addr <= 2'h0;
      end else if (_r_superpage_repl_addr_T_4[1]) begin // @[Mux.scala 47:69]
        r_superpage_repl_addr <= 2'h1;
      end else begin
        r_superpage_repl_addr <= _r_superpage_repl_addr_T_9;
      end
    end
    if (_T_42) begin // @[TLB.scala 359:38]
      if (&r_sectored_repl_addr_valids) begin // @[TLB.scala 407:8]
        r_sectored_repl_addr <= _r_sectored_repl_addr_T_6;
      end else if (_r_sectored_repl_addr_T_8[0]) begin // @[Mux.scala 47:69]
        r_sectored_repl_addr <= 3'h0;
      end else if (_r_sectored_repl_addr_T_8[1]) begin // @[Mux.scala 47:69]
        r_sectored_repl_addr <= 3'h1;
      end else begin
        r_sectored_repl_addr <= _r_sectored_repl_addr_T_21;
      end
    end
    if (_T_42) begin // @[TLB.scala 359:38]
      r_sectored_hit_addr <= state_reg_touch_way_sized; // @[TLB.scala 365:27]
    end
    if (_T_42) begin // @[TLB.scala 359:38]
      r_sectored_hit <= _T_30; // @[TLB.scala 366:22]
    end
    if (_T_23) begin // @[TLB.scala 325:37]
      if (_T_30) begin // @[TLB.scala 326:28]
        state_reg <= _state_reg_T_16; // @[Replacement.scala 162:15]
      end
    end
    if (_T_23) begin // @[TLB.scala 325:37]
      if (_T_37) begin // @[TLB.scala 327:31]
        state_reg_1 <= _state_reg_1_T_6; // @[Replacement.scala 162:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sectored_entries_0_tag = _RAND_0[26:0];
  _RAND_1 = {2{`RANDOM}};
  sectored_entries_0_data_0 = _RAND_1[34:0];
  _RAND_2 = {2{`RANDOM}};
  sectored_entries_0_data_1 = _RAND_2[34:0];
  _RAND_3 = {2{`RANDOM}};
  sectored_entries_0_data_2 = _RAND_3[34:0];
  _RAND_4 = {2{`RANDOM}};
  sectored_entries_0_data_3 = _RAND_4[34:0];
  _RAND_5 = {1{`RANDOM}};
  sectored_entries_0_valid_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  sectored_entries_0_valid_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  sectored_entries_0_valid_2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  sectored_entries_0_valid_3 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  sectored_entries_1_tag = _RAND_9[26:0];
  _RAND_10 = {2{`RANDOM}};
  sectored_entries_1_data_0 = _RAND_10[34:0];
  _RAND_11 = {2{`RANDOM}};
  sectored_entries_1_data_1 = _RAND_11[34:0];
  _RAND_12 = {2{`RANDOM}};
  sectored_entries_1_data_2 = _RAND_12[34:0];
  _RAND_13 = {2{`RANDOM}};
  sectored_entries_1_data_3 = _RAND_13[34:0];
  _RAND_14 = {1{`RANDOM}};
  sectored_entries_1_valid_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  sectored_entries_1_valid_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  sectored_entries_1_valid_2 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  sectored_entries_1_valid_3 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  sectored_entries_2_tag = _RAND_18[26:0];
  _RAND_19 = {2{`RANDOM}};
  sectored_entries_2_data_0 = _RAND_19[34:0];
  _RAND_20 = {2{`RANDOM}};
  sectored_entries_2_data_1 = _RAND_20[34:0];
  _RAND_21 = {2{`RANDOM}};
  sectored_entries_2_data_2 = _RAND_21[34:0];
  _RAND_22 = {2{`RANDOM}};
  sectored_entries_2_data_3 = _RAND_22[34:0];
  _RAND_23 = {1{`RANDOM}};
  sectored_entries_2_valid_0 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  sectored_entries_2_valid_1 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  sectored_entries_2_valid_2 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  sectored_entries_2_valid_3 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  sectored_entries_3_tag = _RAND_27[26:0];
  _RAND_28 = {2{`RANDOM}};
  sectored_entries_3_data_0 = _RAND_28[34:0];
  _RAND_29 = {2{`RANDOM}};
  sectored_entries_3_data_1 = _RAND_29[34:0];
  _RAND_30 = {2{`RANDOM}};
  sectored_entries_3_data_2 = _RAND_30[34:0];
  _RAND_31 = {2{`RANDOM}};
  sectored_entries_3_data_3 = _RAND_31[34:0];
  _RAND_32 = {1{`RANDOM}};
  sectored_entries_3_valid_0 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  sectored_entries_3_valid_1 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  sectored_entries_3_valid_2 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  sectored_entries_3_valid_3 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  sectored_entries_4_tag = _RAND_36[26:0];
  _RAND_37 = {2{`RANDOM}};
  sectored_entries_4_data_0 = _RAND_37[34:0];
  _RAND_38 = {2{`RANDOM}};
  sectored_entries_4_data_1 = _RAND_38[34:0];
  _RAND_39 = {2{`RANDOM}};
  sectored_entries_4_data_2 = _RAND_39[34:0];
  _RAND_40 = {2{`RANDOM}};
  sectored_entries_4_data_3 = _RAND_40[34:0];
  _RAND_41 = {1{`RANDOM}};
  sectored_entries_4_valid_0 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  sectored_entries_4_valid_1 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  sectored_entries_4_valid_2 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  sectored_entries_4_valid_3 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  sectored_entries_5_tag = _RAND_45[26:0];
  _RAND_46 = {2{`RANDOM}};
  sectored_entries_5_data_0 = _RAND_46[34:0];
  _RAND_47 = {2{`RANDOM}};
  sectored_entries_5_data_1 = _RAND_47[34:0];
  _RAND_48 = {2{`RANDOM}};
  sectored_entries_5_data_2 = _RAND_48[34:0];
  _RAND_49 = {2{`RANDOM}};
  sectored_entries_5_data_3 = _RAND_49[34:0];
  _RAND_50 = {1{`RANDOM}};
  sectored_entries_5_valid_0 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  sectored_entries_5_valid_1 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  sectored_entries_5_valid_2 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  sectored_entries_5_valid_3 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  sectored_entries_6_tag = _RAND_54[26:0];
  _RAND_55 = {2{`RANDOM}};
  sectored_entries_6_data_0 = _RAND_55[34:0];
  _RAND_56 = {2{`RANDOM}};
  sectored_entries_6_data_1 = _RAND_56[34:0];
  _RAND_57 = {2{`RANDOM}};
  sectored_entries_6_data_2 = _RAND_57[34:0];
  _RAND_58 = {2{`RANDOM}};
  sectored_entries_6_data_3 = _RAND_58[34:0];
  _RAND_59 = {1{`RANDOM}};
  sectored_entries_6_valid_0 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  sectored_entries_6_valid_1 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  sectored_entries_6_valid_2 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  sectored_entries_6_valid_3 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  sectored_entries_7_tag = _RAND_63[26:0];
  _RAND_64 = {2{`RANDOM}};
  sectored_entries_7_data_0 = _RAND_64[34:0];
  _RAND_65 = {2{`RANDOM}};
  sectored_entries_7_data_1 = _RAND_65[34:0];
  _RAND_66 = {2{`RANDOM}};
  sectored_entries_7_data_2 = _RAND_66[34:0];
  _RAND_67 = {2{`RANDOM}};
  sectored_entries_7_data_3 = _RAND_67[34:0];
  _RAND_68 = {1{`RANDOM}};
  sectored_entries_7_valid_0 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  sectored_entries_7_valid_1 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  sectored_entries_7_valid_2 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  sectored_entries_7_valid_3 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  superpage_entries_0_level = _RAND_72[1:0];
  _RAND_73 = {1{`RANDOM}};
  superpage_entries_0_tag = _RAND_73[26:0];
  _RAND_74 = {2{`RANDOM}};
  superpage_entries_0_data_0 = _RAND_74[34:0];
  _RAND_75 = {1{`RANDOM}};
  superpage_entries_0_valid_0 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  superpage_entries_1_level = _RAND_76[1:0];
  _RAND_77 = {1{`RANDOM}};
  superpage_entries_1_tag = _RAND_77[26:0];
  _RAND_78 = {2{`RANDOM}};
  superpage_entries_1_data_0 = _RAND_78[34:0];
  _RAND_79 = {1{`RANDOM}};
  superpage_entries_1_valid_0 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  superpage_entries_2_level = _RAND_80[1:0];
  _RAND_81 = {1{`RANDOM}};
  superpage_entries_2_tag = _RAND_81[26:0];
  _RAND_82 = {2{`RANDOM}};
  superpage_entries_2_data_0 = _RAND_82[34:0];
  _RAND_83 = {1{`RANDOM}};
  superpage_entries_2_valid_0 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  superpage_entries_3_level = _RAND_84[1:0];
  _RAND_85 = {1{`RANDOM}};
  superpage_entries_3_tag = _RAND_85[26:0];
  _RAND_86 = {2{`RANDOM}};
  superpage_entries_3_data_0 = _RAND_86[34:0];
  _RAND_87 = {1{`RANDOM}};
  superpage_entries_3_valid_0 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  special_entry_level = _RAND_88[1:0];
  _RAND_89 = {1{`RANDOM}};
  special_entry_tag = _RAND_89[26:0];
  _RAND_90 = {2{`RANDOM}};
  special_entry_data_0 = _RAND_90[34:0];
  _RAND_91 = {1{`RANDOM}};
  special_entry_valid_0 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  state = _RAND_92[1:0];
  _RAND_93 = {1{`RANDOM}};
  r_refill_tag = _RAND_93[26:0];
  _RAND_94 = {1{`RANDOM}};
  r_superpage_repl_addr = _RAND_94[1:0];
  _RAND_95 = {1{`RANDOM}};
  r_sectored_repl_addr = _RAND_95[2:0];
  _RAND_96 = {1{`RANDOM}};
  r_sectored_hit_addr = _RAND_96[2:0];
  _RAND_97 = {1{`RANDOM}};
  r_sectored_hit = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  state_reg = _RAND_98[6:0];
  _RAND_99 = {1{`RANDOM}};
  state_reg_1 = _RAND_99[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
