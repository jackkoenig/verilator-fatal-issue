module IntSyncSyncCrossingSink_1(
  input   auto_in_sync_0,
  output  auto_out_0
);
  assign auto_out_0 = auto_in_sync_0; // @[Nodes.scala 1216:84 LazyModule.scala 312:16]
endmodule
