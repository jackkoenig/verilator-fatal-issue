module RecFNToIN_1(
  input  [64:0] io_in,
  input  [2:0]  io_roundingMode,
  input         io_signedOut,
  output [2:0]  io_intExceptionFlags
);
  wire [11:0] rawIn_exp = io_in[63:52]; // @[rawFloatFromRecFN.scala 50:21]
  wire  rawIn_isZero = (rawIn_exp[11:9]) == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  wire  rawIn_isSpecial = (rawIn_exp[11:10]) == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawIn__isNaN = rawIn_isSpecial & (rawIn_exp[9]); // @[rawFloatFromRecFN.scala 55:33]
  wire  rawIn__isInf = rawIn_isSpecial & (~(rawIn_exp[9])); // @[rawFloatFromRecFN.scala 56:33]
  wire  rawIn__sign = io_in[64]; // @[rawFloatFromRecFN.scala 58:25]
  wire [12:0] rawIn__sExp = {1'b0,$signed(rawIn_exp)}; // @[rawFloatFromRecFN.scala 59:27]
  wire  rawIn_rawIn_sig_right_left = ~rawIn_isZero; // @[rawFloatFromRecFN.scala 60:39]
  wire [51:0] rawIn_rawIn_sig_left = io_in[51:0]; // @[rawFloatFromRecFN.scala 60:51]
  wire [53:0] rawIn__sig = {1'h0,rawIn_rawIn_sig_right_left,rawIn_rawIn_sig_left}; // @[Cat.scala 29:58]
  wire  magGeOne = rawIn__sExp[11]; // @[RecFNToIN.scala 58:30]
  wire [10:0] posExp = rawIn__sExp[10:0]; // @[RecFNToIN.scala 59:28]
  wire  magJustBelowOne = (~magGeOne) & (&posExp); // @[RecFNToIN.scala 60:37]
  wire  roundingMode_near_even = io_roundingMode == 3'h0; // @[RecFNToIN.scala 64:53]
  wire  roundingMode_min = io_roundingMode == 3'h2; // @[RecFNToIN.scala 66:53]
  wire  roundingMode_max = io_roundingMode == 3'h3; // @[RecFNToIN.scala 67:53]
  wire  roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RecFNToIN.scala 68:53]
  wire  roundingMode_odd = io_roundingMode == 3'h6; // @[RecFNToIN.scala 69:53]
  wire [51:0] shiftedSig_left = rawIn__sig[51:0]; // @[RecFNToIN.scala 80:32]
  wire [52:0] _shiftedSig_T = {magGeOne,shiftedSig_left}; // @[Cat.scala 29:58]
  wire [4:0] _shiftedSig_T_2 = magGeOne ? rawIn__sExp[4:0] : 5'h0; // @[RecFNToIN.scala 81:16]
  wire [83:0] _GEN_0 = {{31'd0}, _shiftedSig_T}; // @[RecFNToIN.scala 80:50]
  wire [83:0] shiftedSig = _GEN_0 << _shiftedSig_T_2; // @[RecFNToIN.scala 80:50]
  wire [32:0] alignedSig_right = shiftedSig[83:51]; // @[RecFNToIN.scala 86:23]
  wire  alignedSig_left = |(shiftedSig[50:0]); // @[RecFNToIN.scala 86:69]
  wire [33:0] alignedSig = {alignedSig_right,alignedSig_left}; // @[Cat.scala 29:58]
  wire [31:0] unroundedInt = alignedSig[33:2]; // @[RecFNToIN.scala 87:54]
  wire  _common_inexact_T_1 = |(alignedSig[1:0]); // @[RecFNToIN.scala 89:57]
  wire  common_inexact = magGeOne ? |(alignedSig[1:0]) : rawIn_rawIn_sig_right_left; // @[RecFNToIN.scala 89:29]
  wire  _roundIncr_near_even_T_8 = magJustBelowOne & _common_inexact_T_1; // @[RecFNToIN.scala 92:26]
  wire  roundIncr_near_even = (magGeOne & ((&(alignedSig[2:1])) | (&(alignedSig[1:0])))) | _roundIncr_near_even_T_8; // @[RecFNToIN.scala 91:78]
  wire  roundIncr_near_maxMag = (magGeOne & (alignedSig[1])) | magJustBelowOne; // @[RecFNToIN.scala 93:61]
  wire  _roundIncr_T_1 = roundingMode_near_maxMag & roundIncr_near_maxMag; // @[RecFNToIN.scala 96:35]
  wire  _roundIncr_T_2 = (roundingMode_near_even & roundIncr_near_even) | _roundIncr_T_1; // @[RecFNToIN.scala 95:61]
  wire  _roundIncr_T_4 = rawIn__sign & common_inexact; // @[RecFNToIN.scala 98:26]
  wire  _roundIncr_T_5 = (roundingMode_min | roundingMode_odd) & _roundIncr_T_4; // @[RecFNToIN.scala 97:49]
  wire  _roundIncr_T_6 = _roundIncr_T_2 | _roundIncr_T_5; // @[RecFNToIN.scala 96:61]
  wire  _roundIncr_T_9 = roundingMode_max & ((~rawIn__sign) & common_inexact); // @[RecFNToIN.scala 99:27]
  wire  roundIncr = _roundIncr_T_6 | _roundIncr_T_9; // @[RecFNToIN.scala 98:46]
  wire  magGeOne_atOverflowEdge = posExp == 11'h1f; // @[RecFNToIN.scala 107:43]
  wire  roundCarryBut2 = (&(unroundedInt[29:0])) & roundIncr; // @[RecFNToIN.scala 110:61]
  wire  _common_overflow_T_3 = (|(unroundedInt[30:0])) | roundIncr; // @[RecFNToIN.scala 117:64]
  wire  _common_overflow_T_4 = magGeOne_atOverflowEdge & _common_overflow_T_3; // @[RecFNToIN.scala 116:49]
  wire  _common_overflow_T_6 = (posExp == 11'h1e) & roundCarryBut2; // @[RecFNToIN.scala 119:62]
  wire  _common_overflow_T_7 = magGeOne_atOverflowEdge | _common_overflow_T_6; // @[RecFNToIN.scala 118:49]
  wire  _common_overflow_T_8 = rawIn__sign ? _common_overflow_T_4 : _common_overflow_T_7; // @[RecFNToIN.scala 115:24]
  wire  _common_overflow_T_10 = magGeOne_atOverflowEdge & (unroundedInt[30]); // @[RecFNToIN.scala 122:50]
  wire  _common_overflow_T_11 = _common_overflow_T_10 & roundCarryBut2; // @[RecFNToIN.scala 123:57]
  wire  _common_overflow_T_12 = rawIn__sign | _common_overflow_T_11; // @[RecFNToIN.scala 121:32]
  wire  _common_overflow_T_13 = io_signedOut ? _common_overflow_T_8 : _common_overflow_T_12; // @[RecFNToIN.scala 114:20]
  wire  _common_overflow_T_14 = (posExp >= 11'h20) | _common_overflow_T_13; // @[RecFNToIN.scala 113:40]
  wire  _common_overflow_T_17 = ((~io_signedOut) & rawIn__sign) & roundIncr; // @[RecFNToIN.scala 125:41]
  wire  common_overflow = magGeOne ? _common_overflow_T_14 : _common_overflow_T_17; // @[RecFNToIN.scala 112:12]
  wire  invalidExc = rawIn__isNaN | rawIn__isInf; // @[RecFNToIN.scala 130:34]
  wire  _overflow_T = ~invalidExc; // @[RecFNToIN.scala 131:20]
  wire  overflow = (~invalidExc) & common_overflow; // @[RecFNToIN.scala 131:32]
  wire  inexact = (_overflow_T & (~common_overflow)) & common_inexact; // @[RecFNToIN.scala 132:52]
  wire [1:0] io_intExceptionFlags_right = {invalidExc,overflow}; // @[Cat.scala 29:58]
  assign io_intExceptionFlags = {io_intExceptionFlags_right,inexact}; // @[Cat.scala 29:58]
endmodule
